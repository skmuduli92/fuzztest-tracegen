/*verilator coverage_off */

//
// Verific Verilog Description of module oc8051_tb
//

module oc8051_tb (rst, clk, _cvpt_0, _cvpt_1, _cvpt_2, _cvpt_3, 
            _cvpt_4, _cvpt_5, _cvpt_6, _cvpt_7, _cvpt_8, _cvpt_9, 
            _cvpt_10, _cvpt_11, _cvpt_12, _cvpt_13, _cvpt_14, _cvpt_15, 
            _cvpt_16, _cvpt_17, _cvpt_18, _cvpt_19, _cvpt_20, _cvpt_21, 
            _cvpt_22, _cvpt_23, _cvpt_24, _cvpt_25, _cvpt_26, _cvpt_27, 
            _cvpt_28, _cvpt_29, _cvpt_30, _cvpt_31, _cvpt_32, _cvpt_33, 
            _cvpt_34, _cvpt_35, _cvpt_36, _cvpt_37, _cvpt_38, _cvpt_39, 
            _cvpt_40, _cvpt_41, _cvpt_42, _cvpt_43, _cvpt_44, _cvpt_45, 
            _cvpt_46, _cvpt_47, _cvpt_48, _cvpt_49, _cvpt_50, _cvpt_51, 
            _cvpt_52, _cvpt_53, _cvpt_54, _cvpt_55, _cvpt_56, _cvpt_57, 
            _cvpt_58, _cvpt_59, _cvpt_60, _cvpt_61, _cvpt_62, _cvpt_63, 
            _cvpt_64, _cvpt_65, _cvpt_66, _cvpt_67, _cvpt_68, _cvpt_69, 
            _cvpt_70, _cvpt_71, _cvpt_72, _cvpt_73, _cvpt_74, _cvpt_75, 
            _cvpt_76, _cvpt_77, _cvpt_78, _cvpt_79, _cvpt_80, _cvpt_81, 
            _cvpt_82, _cvpt_83, _cvpt_84, _cvpt_85, _cvpt_86, _cvpt_87, 
            _cvpt_88, _cvpt_89, _cvpt_90, _cvpt_91, _cvpt_92, _cvpt_93, 
            _cvpt_94, _cvpt_95, _cvpt_96, _cvpt_97, _cvpt_98, _cvpt_99, 
            _cvpt_100, _cvpt_101, _cvpt_102, _cvpt_103, _cvpt_104, 
            _cvpt_105, _cvpt_106, _cvpt_107, _cvpt_108, _cvpt_109, 
            _cvpt_110, _cvpt_111, _cvpt_112, _cvpt_113, _cvpt_114, 
            _cvpt_115, _cvpt_116, _cvpt_117, _cvpt_118, _cvpt_119, 
            _cvpt_120, _cvpt_121, _cvpt_122, _cvpt_123, _cvpt_124, 
            _cvpt_125, _cvpt_126, _cvpt_127, _cvpt_128, _cvpt_129, 
            _cvpt_130, _cvpt_131, _cvpt_132, _cvpt_133, _cvpt_134, 
            _cvpt_135, _cvpt_136, _cvpt_137, _cvpt_138, _cvpt_139, 
            _cvpt_140, _cvpt_141, _cvpt_142, _cvpt_143, _cvpt_144, 
            _cvpt_145, _cvpt_146, _cvpt_147, _cvpt_148, _cvpt_149, 
            _cvpt_150, _cvpt_151, _cvpt_152, _cvpt_153, _cvpt_154, 
            _cvpt_155, _cvpt_156, _cvpt_157, _cvpt_158, _cvpt_159, 
            _cvpt_160, _cvpt_161, _cvpt_162, _cvpt_163, _cvpt_164, 
            _cvpt_165, _cvpt_166, _cvpt_167, _cvpt_168, _cvpt_169, 
            _cvpt_170, _cvpt_171, _cvpt_172, _cvpt_173, _cvpt_174, 
            _cvpt_175, _cvpt_176, _cvpt_177, _cvpt_178, _cvpt_179, 
            _cvpt_180, _cvpt_181, _cvpt_182, _cvpt_183, _cvpt_184, 
            _cvpt_185, _cvpt_186, _cvpt_187, _cvpt_188, _cvpt_189, 
            _cvpt_190, _cvpt_191, _cvpt_192, _cvpt_193, _cvpt_194, 
            _cvpt_195, _cvpt_196, _cvpt_197, _cvpt_198, _cvpt_199, 
            _cvpt_200, _cvpt_201, _cvpt_202, _cvpt_203, _cvpt_204, 
            _cvpt_205, _cvpt_206, _cvpt_207, _cvpt_208, _cvpt_209, 
            _cvpt_210, _cvpt_211, _cvpt_212, _cvpt_213, _cvpt_214, 
            _cvpt_215, _cvpt_216, _cvpt_217, _cvpt_218, _cvpt_219, 
            _cvpt_220, _cvpt_221, _cvpt_222, _cvpt_223, _cvpt_224, 
            _cvpt_225, _cvpt_226, _cvpt_227, _cvpt_228, _cvpt_229, 
            _cvpt_230, _cvpt_231, _cvpt_232, _cvpt_233, _cvpt_234, 
            _cvpt_235, _cvpt_236, _cvpt_237, _cvpt_238, _cvpt_239, 
            _cvpt_240, _cvpt_241, _cvpt_242, _cvpt_243, _cvpt_244, 
            _cvpt_245, _cvpt_246, _cvpt_247, _cvpt_248, _cvpt_249, 
            _cvpt_250, _cvpt_251, _cvpt_252, _cvpt_253, _cvpt_254, 
            _cvpt_255, _cvpt_256, _cvpt_257, _cvpt_258, _cvpt_259, 
            _cvpt_260, _cvpt_261, _cvpt_262, _cvpt_263, _cvpt_264, 
            _cvpt_265, _cvpt_266, _cvpt_267, _cvpt_268, _cvpt_269, 
            _cvpt_270, _cvpt_271, _cvpt_272, _cvpt_273, _cvpt_274, 
            _cvpt_275, _cvpt_276, _cvpt_277, _cvpt_278, _cvpt_279, 
            _cvpt_280, _cvpt_281, _cvpt_282, _cvpt_283, _cvpt_284, 
            _cvpt_285, _cvpt_286, _cvpt_287, _cvpt_288, _cvpt_289, 
            _cvpt_290, _cvpt_291, _cvpt_292, _cvpt_293, _cvpt_294, 
            _cvpt_295, _cvpt_296, _cvpt_297, _cvpt_298, _cvpt_299, 
            _cvpt_300, _cvpt_301, _cvpt_302, _cvpt_303, _cvpt_304, 
            _cvpt_305, _cvpt_306, _cvpt_307, _cvpt_308, _cvpt_309, 
            _cvpt_310, _cvpt_311, _cvpt_312, _cvpt_313, _cvpt_314, 
            _cvpt_315, _cvpt_316, _cvpt_317, _cvpt_318, _cvpt_319, 
            _cvpt_320, _cvpt_321, _cvpt_322, _cvpt_323, _cvpt_324, 
            _cvpt_325, _cvpt_326, _cvpt_327, _cvpt_328, _cvpt_329, 
            _cvpt_330, _cvpt_331, _cvpt_332, _cvpt_333, _cvpt_334, 
            _cvpt_335, _cvpt_336, _cvpt_337, _cvpt_338, _cvpt_339, 
            _cvpt_340, _cvpt_341, _cvpt_342, _cvpt_343, _cvpt_344, 
            _cvpt_345, _cvpt_346, _cvpt_347, _cvpt_348, _cvpt_349, 
            _cvpt_350, _cvpt_351, _cvpt_352, _cvpt_353, _cvpt_354, 
            _cvpt_355, _cvpt_356, _cvpt_357, _cvpt_358, _cvpt_359, 
            _cvpt_360, _cvpt_361, _cvpt_362, _cvpt_363, _cvpt_364, 
            _cvpt_365, _cvpt_366, _cvpt_367, _cvpt_368, _cvpt_369, 
            _cvpt_370, _cvpt_371, _cvpt_372, _cvpt_373, _cvpt_374, 
            _cvpt_375, _cvpt_376, _cvpt_377, _cvpt_378, _cvpt_379, 
            _cvpt_380, _cvpt_381, _cvpt_382, _cvpt_383, _cvpt_384, 
            _cvpt_385, _cvpt_386, _cvpt_387, _cvpt_388, _cvpt_389, 
            _cvpt_390, _cvpt_391, _cvpt_392, _cvpt_393, _cvpt_394, 
            _cvpt_395, _cvpt_396, _cvpt_397, _cvpt_398, _cvpt_399, 
            _cvpt_400, _cvpt_401, _cvpt_402, _cvpt_403, _cvpt_404, 
            _cvpt_405, _cvpt_406, _cvpt_407, _cvpt_408, _cvpt_409, 
            _cvpt_410, _cvpt_411, _cvpt_412, _cvpt_413, _cvpt_414, 
            _cvpt_415, _cvpt_416, _cvpt_417, _cvpt_418, _cvpt_419, 
            _cvpt_420, _cvpt_421, _cvpt_422, _cvpt_423, _cvpt_424, 
            _cvpt_425, _cvpt_426, _cvpt_427, _cvpt_428, _cvpt_429, 
            _cvpt_430, _cvpt_431, _cvpt_432, _cvpt_433, _cvpt_434, 
            _cvpt_435, _cvpt_436, _cvpt_437, _cvpt_438, _cvpt_439, 
            _cvpt_440, _cvpt_441, _cvpt_442, _cvpt_443, _cvpt_444, 
            _cvpt_445, _cvpt_446, _cvpt_447, _cvpt_448, _cvpt_449, 
            _cvpt_450, _cvpt_451, _cvpt_452, _cvpt_453, _cvpt_454, 
            _cvpt_455, _cvpt_456, _cvpt_457, _cvpt_458, _cvpt_459, 
            _cvpt_460, _cvpt_461, _cvpt_462, _cvpt_463, _cvpt_464, 
            _cvpt_465, _cvpt_466, _cvpt_467, _cvpt_468, _cvpt_469, 
            _cvpt_470, _cvpt_471, _cvpt_472, _cvpt_473, _cvpt_474, 
            _cvpt_475, _cvpt_476, _cvpt_477, _cvpt_478, _cvpt_479, 
            _cvpt_480, _cvpt_481, _cvpt_482, _cvpt_483, _cvpt_484, 
            _cvpt_485, _cvpt_486, _cvpt_487, _cvpt_488, _cvpt_489, 
            _cvpt_490, _cvpt_491, _cvpt_492, _cvpt_493, _cvpt_494, 
            _cvpt_495, _cvpt_496, _cvpt_497, _cvpt_498, _cvpt_499, 
            _cvpt_500, _cvpt_501, _cvpt_502, _cvpt_503, _cvpt_504, 
            _cvpt_505, _cvpt_506, _cvpt_507, _cvpt_508, _cvpt_509, 
            _cvpt_510, _cvpt_511, _cvpt_512, _cvpt_513, _cvpt_514, 
            _cvpt_515, _cvpt_516, _cvpt_517, _cvpt_518, _cvpt_519, 
            _cvpt_520, _cvpt_521, _cvpt_522, _cvpt_523, _cvpt_524, 
            _cvpt_525, _cvpt_526, _cvpt_527, _cvpt_528, _cvpt_529, 
            _cvpt_530, _cvpt_531, _cvpt_532, _cvpt_533, _cvpt_534, 
            _cvpt_535, _cvpt_536, _cvpt_537, _cvpt_538, _cvpt_539, 
            _cvpt_540, _cvpt_541, _cvpt_542, _cvpt_543, _cvpt_544, 
            _cvpt_545, _cvpt_546, _cvpt_547, _cvpt_548, _cvpt_549, 
            _cvpt_550, _cvpt_551, _cvpt_552, _cvpt_553, _cvpt_554, 
            _cvpt_555, _cvpt_556, _cvpt_557, _cvpt_558, _cvpt_559, 
            _cvpt_560, _cvpt_561, _cvpt_562, _cvpt_563, _cvpt_564, 
            _cvpt_565, _cvpt_566, _cvpt_567, _cvpt_568, _cvpt_569, 
            _cvpt_570, _cvpt_571, _cvpt_572, _cvpt_573, _cvpt_574, 
            _cvpt_575, _cvpt_576, _cvpt_577, _cvpt_578, _cvpt_579, 
            _cvpt_580, _cvpt_581, _cvpt_582, _cvpt_583, _cvpt_584, 
            _cvpt_585, _cvpt_586, _cvpt_587, _cvpt_588, _cvpt_589, 
            _cvpt_590, _cvpt_591, _cvpt_592, _cvpt_593, _cvpt_594, 
            _cvpt_595, _cvpt_596, _cvpt_597, _cvpt_598, _cvpt_599, 
            _cvpt_600, _cvpt_601, _cvpt_602, _cvpt_603, _cvpt_604, 
            _cvpt_605, _cvpt_606, _cvpt_607, _cvpt_608, _cvpt_609, 
            _cvpt_610, _cvpt_611, _cvpt_612, _cvpt_613, _cvpt_614, 
            _cvpt_615, _cvpt_616, _cvpt_617, _cvpt_618, _cvpt_619, 
            _cvpt_620, _cvpt_621, _cvpt_622, _cvpt_623, _cvpt_624, 
            _cvpt_625, _cvpt_626, _cvpt_627, _cvpt_628, _cvpt_629, 
            _cvpt_630, _cvpt_631, _cvpt_632, _cvpt_633, _cvpt_634, 
            _cvpt_635, _cvpt_636, _cvpt_637, _cvpt_638, _cvpt_639, 
            _cvpt_640, _cvpt_641, _cvpt_642, _cvpt_643, _cvpt_644, 
            _cvpt_645, _cvpt_646, _cvpt_647, _cvpt_648, _cvpt_649, 
            _cvpt_650, _cvpt_651, _cvpt_652, _cvpt_653, _cvpt_654, 
            _cvpt_655, _cvpt_656, _cvpt_657, _cvpt_658, _cvpt_659, 
            _cvpt_660, _cvpt_661, _cvpt_662, _cvpt_663, _cvpt_664, 
            _cvpt_665, _cvpt_666, _cvpt_667, _cvpt_668, _cvpt_669, 
            _cvpt_670, _cvpt_671, _cvpt_672, _cvpt_673, _cvpt_674, 
            _cvpt_675, _cvpt_676, _cvpt_677, _cvpt_678, _cvpt_679, 
            _cvpt_680, _cvpt_681, _cvpt_682, _cvpt_683, _cvpt_684, 
            _cvpt_685, _cvpt_686, _cvpt_687, _cvpt_688, _cvpt_689, 
            _cvpt_690, _cvpt_691, _cvpt_692, _cvpt_693, _cvpt_694, 
            _cvpt_695, _cvpt_696, _cvpt_697, _cvpt_698, _cvpt_699, 
            _cvpt_700, _cvpt_701, _cvpt_702, _cvpt_703, _cvpt_704, 
            _cvpt_705, _cvpt_706, _cvpt_707, _cvpt_708, _cvpt_709, 
            _cvpt_710, _cvpt_711, _cvpt_712, _cvpt_713, _cvpt_714, 
            _cvpt_715, _cvpt_716, _cvpt_717, _cvpt_718, _cvpt_719, 
            _cvpt_720, _cvpt_721, _cvpt_722, _cvpt_723, _cvpt_724, 
            _cvpt_725, _cvpt_726, _cvpt_727, _cvpt_728, _cvpt_729, 
            _cvpt_730, _cvpt_731, _cvpt_732, _cvpt_733, _cvpt_734, 
            _cvpt_735, _cvpt_736, _cvpt_737, _cvpt_738, _cvpt_739, 
            _cvpt_740, _cvpt_741, _cvpt_742, _cvpt_743, _cvpt_744, 
            _cvpt_745, _cvpt_746, _cvpt_747, _cvpt_748, _cvpt_749, 
            _cvpt_750, _cvpt_751, _cvpt_752, _cvpt_753, _cvpt_754, 
            _cvpt_755, _cvpt_756, _cvpt_757, _cvpt_758, _cvpt_759, 
            _cvpt_760, _cvpt_761, _cvpt_762, _cvpt_763, _cvpt_764, 
            _cvpt_765, _cvpt_766, _cvpt_767, _cvpt_768, _cvpt_769, 
            _cvpt_770, _cvpt_771, _cvpt_772, _cvpt_773, _cvpt_774, 
            _cvpt_775, _cvpt_776, _cvpt_777, _cvpt_778, _cvpt_779, 
            _cvpt_780, _cvpt_781, _cvpt_782, _cvpt_783, _cvpt_784, 
            _cvpt_785, _cvpt_786, _cvpt_787, _cvpt_788, _cvpt_789, 
            _cvpt_790, _cvpt_791, _cvpt_792, _cvpt_793, _cvpt_794, 
            _cvpt_795, _cvpt_796, _cvpt_797, _cvpt_798, _cvpt_799, 
            _cvpt_800, _cvpt_801, _cvpt_802, _cvpt_803, _cvpt_804, 
            _cvpt_805, _cvpt_806, _cvpt_807, _cvpt_808, _cvpt_809, 
            _cvpt_810, _cvpt_811, _cvpt_812, _cvpt_813, _cvpt_814, 
            _cvpt_815, _cvpt_816, _cvpt_817, _cvpt_818, _cvpt_819, 
            _cvpt_820, _cvpt_821, _cvpt_822, _cvpt_823, _cvpt_824, 
            _cvpt_825, _cvpt_826, _cvpt_827, _cvpt_828, _cvpt_829, 
            _cvpt_830, _cvpt_831, _cvpt_832, _cvpt_833, _cvpt_834, 
            _cvpt_835, _cvpt_836, _cvpt_837, _cvpt_838, _cvpt_839, 
            _cvpt_840, _cvpt_841, _cvpt_842, _cvpt_843, _cvpt_844, 
            _cvpt_845, _cvpt_846, _cvpt_847, _cvpt_848, _cvpt_849, 
            _cvpt_850, _cvpt_851, _cvpt_852, _cvpt_853, _cvpt_854, 
            _cvpt_855, _cvpt_856, _cvpt_857, _cvpt_858, _cvpt_859, 
            _cvpt_860, _cvpt_861, _cvpt_862, _cvpt_863, _cvpt_864, 
            _cvpt_865, _cvpt_866, _cvpt_867, _cvpt_868, _cvpt_869, 
            _cvpt_870, _cvpt_871, _cvpt_872, _cvpt_873, _cvpt_874, 
            _cvpt_875, _cvpt_876, _cvpt_877, _cvpt_878, _cvpt_879, 
            _cvpt_880, _cvpt_881, _cvpt_882, _cvpt_883, _cvpt_884, 
            _cvpt_885, _cvpt_886, _cvpt_887, _cvpt_888, _cvpt_889, 
            _cvpt_890, _cvpt_891, _cvpt_892, _cvpt_893, _cvpt_894, 
            _cvpt_895, _cvpt_896, _cvpt_897, _cvpt_898, _cvpt_899, 
            _cvpt_900, _cvpt_901, _cvpt_902, _cvpt_903, _cvpt_904, 
            _cvpt_905, _cvpt_906, _cvpt_907, _cvpt_908, _cvpt_909, 
            _cvpt_910, _cvpt_911, _cvpt_912, _cvpt_913, _cvpt_914, 
            _cvpt_915, _cvpt_916, _cvpt_917, _cvpt_918, _cvpt_919, 
            _cvpt_920, _cvpt_921, _cvpt_922, _cvpt_923, _cvpt_924, 
            _cvpt_925, _cvpt_926, _cvpt_927, _cvpt_928, _cvpt_929, 
            _cvpt_930, _cvpt_931, _cvpt_932, _cvpt_933, _cvpt_934, 
            _cvpt_935, _cvpt_936, _cvpt_937, _cvpt_938, _cvpt_939, 
            _cvpt_940, _cvpt_941, _cvpt_942, _cvpt_943, _cvpt_944, 
            _cvpt_945, _cvpt_946, _cvpt_947, _cvpt_948, _cvpt_949, 
            _cvpt_950, _cvpt_951, _cvpt_952, _cvpt_953, _cvpt_954, 
            _cvpt_955, _cvpt_956, _cvpt_957, _cvpt_958, _cvpt_959, 
            _cvpt_960, _cvpt_961, _cvpt_962, _cvpt_963, _cvpt_964, 
            _cvpt_965, _cvpt_966, _cvpt_967, _cvpt_968, _cvpt_969, 
            _cvpt_970, _cvpt_971, _cvpt_972, _cvpt_973, _cvpt_974, 
            _cvpt_975, _cvpt_976, _cvpt_977, _cvpt_978, _cvpt_979, 
            _cvpt_980, _cvpt_981, _cvpt_982, _cvpt_983, _cvpt_984, 
            _cvpt_985, _cvpt_986, _cvpt_987, _cvpt_988, _cvpt_989, 
            _cvpt_990, _cvpt_991, _cvpt_992, _cvpt_993, _cvpt_994, 
            _cvpt_995, _cvpt_996, _cvpt_997, _cvpt_998, _cvpt_999, 
            _cvpt_1000, _cvpt_1001, _cvpt_1002, _cvpt_1003, _cvpt_1004, 
            _cvpt_1005, _cvpt_1006, _cvpt_1007, _cvpt_1008, _cvpt_1009, 
            _cvpt_1010, _cvpt_1011, _cvpt_1012, _cvpt_1013, _cvpt_1014, 
            _cvpt_1015, _cvpt_1016, _cvpt_1017, _cvpt_1018, _cvpt_1019, 
            _cvpt_1020, _cvpt_1021, _cvpt_1022, _cvpt_1023, _cvpt_1024, 
            _cvpt_1025, _cvpt_1026, _cvpt_1027, _cvpt_1028, _cvpt_1029, 
            _cvpt_1030, _cvpt_1031, _cvpt_1032, _cvpt_1033, _cvpt_1034, 
            _cvpt_1035, _cvpt_1036, _cvpt_1037, _cvpt_1038, _cvpt_1039, 
            _cvpt_1040, _cvpt_1041, _cvpt_1042, _cvpt_1043, _cvpt_1044, 
            _cvpt_1045, _cvpt_1046, _cvpt_1047, _cvpt_1048, _cvpt_1049, 
            _cvpt_1050, _cvpt_1051, _cvpt_1052, _cvpt_1053, _cvpt_1054, 
            _cvpt_1055, _cvpt_1056, _cvpt_1057, _cvpt_1058, _cvpt_1059, 
            _cvpt_1060, _cvpt_1061, _cvpt_1062, _cvpt_1063, _cvpt_1064, 
            _cvpt_1065, _cvpt_1066, _cvpt_1067, _cvpt_1068, _cvpt_1069, 
            _cvpt_1070, _cvpt_1071, _cvpt_1072, _cvpt_1073, _cvpt_1074, 
            _cvpt_1075, _cvpt_1076, _cvpt_1077, _cvpt_1078, _cvpt_1079, 
            _cvpt_1080, _cvpt_1081, _cvpt_1082, _cvpt_1083, _cvpt_1084, 
            _cvpt_1085, _cvpt_1086, _cvpt_1087, _cvpt_1088, _cvpt_1089, 
            _cvpt_1090, _cvpt_1091, _cvpt_1092, _cvpt_1093, _cvpt_1094, 
            _cvpt_1095, _cvpt_1096, _cvpt_1097, _cvpt_1098, _cvpt_1099, 
            _cvpt_1100, _cvpt_1101, _cvpt_1102, _cvpt_1103, _cvpt_1104, 
            _cvpt_1105, _cvpt_1106, _cvpt_1107, _cvpt_1108, _cvpt_1109, 
            _cvpt_1110, _cvpt_1111, _cvpt_1112, _cvpt_1113, _cvpt_1114, 
            _cvpt_1115, _cvpt_1116, _cvpt_1117, _cvpt_1118, _cvpt_1119, 
            _cvpt_1120, _cvpt_1121, _cvpt_1122, _cvpt_1123, _cvpt_1124, 
            _cvpt_1125, _cvpt_1126, _cvpt_1127, _cvpt_1128, _cvpt_1129, 
            _cvpt_1130, _cvpt_1131, _cvpt_1132, _cvpt_1133, _cvpt_1134, 
            _cvpt_1135, _cvpt_1136, _cvpt_1137, _cvpt_1138, _cvpt_1139, 
            _cvpt_1140, _cvpt_1141, _cvpt_1142, _cvpt_1143, _cvpt_1144, 
            _cvpt_1145, _cvpt_1146, _cvpt_1147, _cvpt_1148, _cvpt_1149, 
            _cvpt_1150, _cvpt_1151, _cvpt_1152, _cvpt_1153, _cvpt_1154, 
            _cvpt_1155, _cvpt_1156, _cvpt_1157, _cvpt_1158, _cvpt_1159, 
            _cvpt_1160, _cvpt_1161, _cvpt_1162, _cvpt_1163, _cvpt_1164, 
            _cvpt_1165, _cvpt_1166, _cvpt_1167, _cvpt_1168, _cvpt_1169, 
            _cvpt_1170, _cvpt_1171, _cvpt_1172, _cvpt_1173, _cvpt_1174, 
            _cvpt_1175, _cvpt_1176, _cvpt_1177, _cvpt_1178, _cvpt_1179, 
            _cvpt_1180, _cvpt_1181, _cvpt_1182, _cvpt_1183, _cvpt_1184, 
            _cvpt_1185, _cvpt_1186, _cvpt_1187, _cvpt_1188, _cvpt_1189, 
            _cvpt_1190, _cvpt_1191, _cvpt_1192, _cvpt_1193, _cvpt_1194, 
            _cvpt_1195, _cvpt_1196, _cvpt_1197, _cvpt_1198, _cvpt_1199, 
            _cvpt_1200, _cvpt_1201, _cvpt_1202, _cvpt_1203, _cvpt_1204, 
            _cvpt_1205, _cvpt_1206, _cvpt_1207, _cvpt_1208, _cvpt_1209, 
            _cvpt_1210, _cvpt_1211, _cvpt_1212, _cvpt_1213, _cvpt_1214, 
            _cvpt_1215, _cvpt_1216, _cvpt_1217, _cvpt_1218, _cvpt_1219, 
            _cvpt_1220, _cvpt_1221, _cvpt_1222, _cvpt_1223, _cvpt_1224, 
            _cvpt_1225, _cvpt_1226, _cvpt_1227, _cvpt_1228, _cvpt_1229, 
            _cvpt_1230, _cvpt_1231, _cvpt_1232, _cvpt_1233, _cvpt_1234, 
            _cvpt_1235, _cvpt_1236, _cvpt_1237, _cvpt_1238, _cvpt_1239, 
            _cvpt_1240, _cvpt_1241, _cvpt_1242, _cvpt_1243, _cvpt_1244, 
            _cvpt_1245, _cvpt_1246, _cvpt_1247, _cvpt_1248, _cvpt_1249, 
            _cvpt_1250, _cvpt_1251, _cvpt_1252, _cvpt_1253, _cvpt_1254, 
            _cvpt_1255, _cvpt_1256, _cvpt_1257, _cvpt_1258, _cvpt_1259, 
            _cvpt_1260, _cvpt_1261, _cvpt_1262, _cvpt_1263, _cvpt_1264, 
            _cvpt_1265, _cvpt_1266, _cvpt_1267, _cvpt_1268, _cvpt_1269, 
            _cvpt_1270, _cvpt_1271, _cvpt_1272, _cvpt_1273, _cvpt_1274, 
            _cvpt_1275, _cvpt_1276, _cvpt_1277, _cvpt_1278, _cvpt_1279, 
            _cvpt_1280, _cvpt_1281, _cvpt_1282, _cvpt_1283, _cvpt_1284, 
            _cvpt_1285, _cvpt_1286, _cvpt_1287, _cvpt_1288, _cvpt_1289, 
            _cvpt_1290, _cvpt_1291, _cvpt_1292, _cvpt_1293, _cvpt_1294, 
            _cvpt_1295, _cvpt_1296, _cvpt_1297, _cvpt_1298, _cvpt_1299, 
            _cvpt_1300, _cvpt_1301, _cvpt_1302, _cvpt_1303, _cvpt_1304, 
            _cvpt_1305, _cvpt_1306, _cvpt_1307, _cvpt_1308, _cvpt_1309, 
            _cvpt_1310, _cvpt_1311, _cvpt_1312, _cvpt_1313, _cvpt_1314, 
            _cvpt_1315, _cvpt_1316, _cvpt_1317, _cvpt_1318, _cvpt_1319, 
            _cvpt_1320, _cvpt_1321, _cvpt_1322, _cvpt_1323, _cvpt_1324, 
            _cvpt_1325, _cvpt_1326, _cvpt_1327, _cvpt_1328, _cvpt_1329, 
            _cvpt_1330, _cvpt_1331, _cvpt_1332, _cvpt_1333, _cvpt_1334, 
            _cvpt_1335, _cvpt_1336, _cvpt_1337, _cvpt_1338, _cvpt_1339, 
            _cvpt_1340, _cvpt_1341, _cvpt_1342, _cvpt_1343, _cvpt_1344, 
            _cvpt_1345, _cvpt_1346, _cvpt_1347, _cvpt_1348, _cvpt_1349, 
            _cvpt_1350, _cvpt_1351, _cvpt_1352, _cvpt_1353, _cvpt_1354, 
            _cvpt_1355, _cvpt_1356, _cvpt_1357, _cvpt_1358, _cvpt_1359, 
            _cvpt_1360, _cvpt_1361, _cvpt_1362, _cvpt_1363, _cvpt_1364, 
            _cvpt_1365, _cvpt_1366, _cvpt_1367, _cvpt_1368, _cvpt_1369, 
            _cvpt_1370, _cvpt_1371, _cvpt_1372, _cvpt_1373, _cvpt_1374, 
            _cvpt_1375, _cvpt_1376, _cvpt_1377, _cvpt_1378, _cvpt_1379, 
            _cvpt_1380, _cvpt_1381, _cvpt_1382, _cvpt_1383, _cvpt_1384, 
            _cvpt_1385, _cvpt_1386, _cvpt_1387, _cvpt_1388, _cvpt_1389, 
            _cvpt_1390, _cvpt_1391, _cvpt_1392, _cvpt_1393, _cvpt_1394, 
            _cvpt_1395, _cvpt_1396, _cvpt_1397, _cvpt_1398, _cvpt_1399, 
            _cvpt_1400, _cvpt_1401, _cvpt_1402, _cvpt_1403, _cvpt_1404, 
            _cvpt_1405, _cvpt_1406, _cvpt_1407, _cvpt_1408, _cvpt_1409, 
            _cvpt_1410, _cvpt_1411, _cvpt_1412, _cvpt_1413, _cvpt_1414, 
            _cvpt_1415, _cvpt_1416, _cvpt_1417, _cvpt_1418, _cvpt_1419, 
            _cvpt_1420, _cvpt_1421, _cvpt_1422, _cvpt_1423, _cvpt_1424, 
            _cvpt_1425, _cvpt_1426, _cvpt_1427, _cvpt_1428, _cvpt_1429, 
            _cvpt_1430, _cvpt_1431, _cvpt_1432, _cvpt_1433, _cvpt_1434, 
            _cvpt_1435, _cvpt_1436, _cvpt_1437, _cvpt_1438, _cvpt_1439, 
            _cvpt_1440, _cvpt_1441, _cvpt_1442, _cvpt_1443, _cvpt_1444, 
            _cvpt_1445, _cvpt_1446, _cvpt_1447, _cvpt_1448, _cvpt_1449, 
            _cvpt_1450, _cvpt_1451, _cvpt_1452, _cvpt_1453, _cvpt_1454, 
            _cvpt_1455, _cvpt_1456, _cvpt_1457, _cvpt_1458, _cvpt_1459, 
            _cvpt_1460, _cvpt_1461, _cvpt_1462, _cvpt_1463, _cvpt_1464, 
            _cvpt_1465, _cvpt_1466, _cvpt_1467, _cvpt_1468, _cvpt_1469, 
            _cvpt_1470, _cvpt_1471, _cvpt_1472, _cvpt_1473, _cvpt_1474, 
            _cvpt_1475, _cvpt_1476, _cvpt_1477, _cvpt_1478, _cvpt_1479, 
            _cvpt_1480, _cvpt_1481, _cvpt_1482, _cvpt_1483, _cvpt_1484, 
            _cvpt_1485, _cvpt_1486, _cvpt_1487, _cvpt_1488, _cvpt_1489, 
            _cvpt_1490, _cvpt_1491, _cvpt_1492, _cvpt_1493, _cvpt_1494, 
            _cvpt_1495, _cvpt_1496, _cvpt_1497, _cvpt_1498, _cvpt_1499, 
            _cvpt_1500, _cvpt_1501, _cvpt_1502, _cvpt_1503, _cvpt_1504, 
            _cvpt_1505, _cvpt_1506, _cvpt_1507, _cvpt_1508, _cvpt_1509, 
            _cvpt_1510, _cvpt_1511, _cvpt_1512, _cvpt_1513, _cvpt_1514, 
            _cvpt_1515, _cvpt_1516, _cvpt_1517, _cvpt_1518, _cvpt_1519, 
            _cvpt_1520, _cvpt_1521, _cvpt_1522, _cvpt_1523, _cvpt_1524, 
            _cvpt_1525, _cvpt_1526, _cvpt_1527, _cvpt_1528, _cvpt_1529, 
            _cvpt_1530, _cvpt_1531, _cvpt_1532, _cvpt_1533, _cvpt_1534, 
            _cvpt_1535, _cvpt_1536, _cvpt_1537, _cvpt_1538, _cvpt_1539, 
            _cvpt_1540, _cvpt_1541, _cvpt_1542, _cvpt_1543, _cvpt_1544, 
            _cvpt_1545, _cvpt_1546, _cvpt_1547, _cvpt_1548, _cvpt_1549, 
            _cvpt_1550, _cvpt_1551, _cvpt_1552, _cvpt_1553, _cvpt_1554, 
            _cvpt_1555, _cvpt_1556, _cvpt_1557, _cvpt_1558, _cvpt_1559, 
            _cvpt_1560, _cvpt_1561, _cvpt_1562, _cvpt_1563, _cvpt_1564, 
            _cvpt_1565, _cvpt_1566, _cvpt_1567, _cvpt_1568, _cvpt_1569, 
            _cvpt_1570, _cvpt_1571, _cvpt_1572, _cvpt_1573, _cvpt_1574, 
            _cvpt_1575, _cvpt_1576, _cvpt_1577, _cvpt_1578, _cvpt_1579, 
            _cvpt_1580, _cvpt_1581, _cvpt_1582, _cvpt_1583, _cvpt_1584, 
            _cvpt_1585, _cvpt_1586, _cvpt_1587, _cvpt_1588, _cvpt_1589, 
            _cvpt_1590, _cvpt_1591, _cvpt_1592, _cvpt_1593, _cvpt_1594, 
            _cvpt_1595, _cvpt_1596, _cvpt_1597, _cvpt_1598, _cvpt_1599, 
            _cvpt_1600, _cvpt_1601, _cvpt_1602, _cvpt_1603, _cvpt_1604, 
            _cvpt_1605, _cvpt_1606, _cvpt_1607, _cvpt_1608, _cvpt_1609, 
            _cvpt_1610, _cvpt_1611, _cvpt_1612, _cvpt_1613, _cvpt_1614, 
            _cvpt_1615, _cvpt_1616, _cvpt_1617, _cvpt_1618, _cvpt_1619, 
            _cvpt_1620, _cvpt_1621, _cvpt_1622, _cvpt_1623, _cvpt_1624, 
            _cvpt_1625, _cvpt_1626, _cvpt_1627, _cvpt_1628, _cvpt_1629, 
            _cvpt_1630, _cvpt_1631, _cvpt_1632, _cvpt_1633, _cvpt_1634, 
            _cvpt_1635, _cvpt_1636, _cvpt_1637, _cvpt_1638, _cvpt_1639, 
            _cvpt_1640, _cvpt_1641, _cvpt_1642, _cvpt_1643, _cvpt_1644, 
            _cvpt_1645, _cvpt_1646, _cvpt_1647, _cvpt_1648, _cvpt_1649, 
            _cvpt_1650, _cvpt_1651, _cvpt_1652, _cvpt_1653, _cvpt_1654, 
            _cvpt_1655, _cvpt_1656, _cvpt_1657, _cvpt_1658, _cvpt_1659, 
            _cvpt_1660, _cvpt_1661, _cvpt_1662, _cvpt_1663, _cvpt_1664, 
            _cvpt_1665, _cvpt_1666, _cvpt_1667, _cvpt_1668, _cvpt_1669, 
            _cvpt_1670, _cvpt_1671, _cvpt_1672, _cvpt_1673, _cvpt_1674, 
            _cvpt_1675, _cvpt_1676, _cvpt_1677, _cvpt_1678, _cvpt_1679, 
            _cvpt_1680, _cvpt_1681, _cvpt_1682, _cvpt_1683, _cvpt_1684, 
            _cvpt_1685, _cvpt_1686, _cvpt_1687, _cvpt_1688, _cvpt_1689, 
            _cvpt_1690, _cvpt_1691, _cvpt_1692, _cvpt_1693, _cvpt_1694, 
            _cvpt_1695, _cvpt_1696, _cvpt_1697, _cvpt_1698, _cvpt_1699, 
            _cvpt_1700, _cvpt_1701, _cvpt_1702, _cvpt_1703, _cvpt_1704, 
            _cvpt_1705, _cvpt_1706, _cvpt_1707, _cvpt_1708, _cvpt_1709, 
            _cvpt_1710, _cvpt_1711, _cvpt_1712, _cvpt_1713, _cvpt_1714, 
            _cvpt_1715, _cvpt_1716, _cvpt_1717, _cvpt_1718, _cvpt_1719, 
            _cvpt_1720, _cvpt_1721, _cvpt_1722, _cvpt_1723, _cvpt_1724, 
            _cvpt_1725, _cvpt_1726, _cvpt_1727, _cvpt_1728, _cvpt_1729, 
            _cvpt_1730, _cvpt_1731, _cvpt_1732, _cvpt_1733, _cvpt_1734, 
            _cvpt_1735, _cvpt_1736, _cvpt_1737, _cvpt_1738, _cvpt_1739, 
            _cvpt_1740, _cvpt_1741, _cvpt_1742, _cvpt_1743, _cvpt_1744, 
            _cvpt_1745, _cvpt_1746, _cvpt_1747, _cvpt_1748, _cvpt_1749, 
            _cvpt_1750, _cvpt_1751, _cvpt_1752, _cvpt_1753, _cvpt_1754, 
            _cvpt_1755, _cvpt_1756, _cvpt_1757, _cvpt_1758, _cvpt_1759, 
            _cvpt_1760, _cvpt_1761, _cvpt_1762, _cvpt_1763, _cvpt_1764, 
            _cvpt_1765, _cvpt_1766, _cvpt_1767, _cvpt_1768, _cvpt_1769, 
            _cvpt_1770, _cvpt_1771, _cvpt_1772, _cvpt_1773, _cvpt_1774, 
            _cvpt_1775, _cvpt_1776, _cvpt_1777, _cvpt_1778, _cvpt_1779, 
            _cvpt_1780, _cvpt_1781, _cvpt_1782, _cvpt_1783, _cvpt_1784, 
            _cvpt_1785, _cvpt_1786, _cvpt_1787, _cvpt_1788, _cvpt_1789, 
            _cvpt_1790, _cvpt_1791, _cvpt_1792, _cvpt_1793, _cvpt_1794, 
            _cvpt_1795, _cvpt_1796, _cvpt_1797, _cvpt_1798, _cvpt_1799, 
            _cvpt_1800, _cvpt_1801, _cvpt_1802, _cvpt_1803, _cvpt_1804, 
            _cvpt_1805, _cvpt_1806, _cvpt_1807, _cvpt_1808, _cvpt_1809, 
            _cvpt_1810, _cvpt_1811, _cvpt_1812, _cvpt_1813, _cvpt_1814, 
            _cvpt_1815, _cvpt_1816, _cvpt_1817, _cvpt_1818, _cvpt_1819, 
            _cvpt_1820, _cvpt_1821, _cvpt_1822, _cvpt_1823, _cvpt_1824, 
            _cvpt_1825, _cvpt_1826, _cvpt_1827, _cvpt_1828, _cvpt_1829, 
            _cvpt_1830, _cvpt_1831, _cvpt_1832, _cvpt_1833, _cvpt_1834, 
            _cvpt_1835, _cvpt_1836, _cvpt_1837, _cvpt_1838, _cvpt_1839, 
            _cvpt_1840, _cvpt_1841, _cvpt_1842, _cvpt_1843, _cvpt_1844, 
            _cvpt_1845, _cvpt_1846, _cvpt_1847, _cvpt_1848, _cvpt_1849, 
            _cvpt_1850, _cvpt_1851, _cvpt_1852, _cvpt_1853, _cvpt_1854, 
            _cvpt_1855, _cvpt_1856, _cvpt_1857, _cvpt_1858, _cvpt_1859, 
            _cvpt_1860, _cvpt_1861, _cvpt_1862, _cvpt_1863, _cvpt_1864, 
            _cvpt_1865, _cvpt_1866, _cvpt_1867, _cvpt_1868, _cvpt_1869, 
            _cvpt_1870, _cvpt_1871, _cvpt_1872, _cvpt_1873, _cvpt_1874, 
            _cvpt_1875, _cvpt_1876, _cvpt_1877, _cvpt_1878, _cvpt_1879, 
            _cvpt_1880, _cvpt_1881, _cvpt_1882, _cvpt_1883, _cvpt_1884, 
            _cvpt_1885, _cvpt_1886, _cvpt_1887, _cvpt_1888, _cvpt_1889, 
            _cvpt_1890, _cvpt_1891, _cvpt_1892, _cvpt_1893, _cvpt_1894, 
            _cvpt_1895, _cvpt_1896, _cvpt_1897, _cvpt_1898, _cvpt_1899, 
            _cvpt_1900, _cvpt_1901, _cvpt_1902, _cvpt_1903, _cvpt_1904, 
            _cvpt_1905, _cvpt_1906, _cvpt_1907, _cvpt_1908, _cvpt_1909, 
            _cvpt_1910, _cvpt_1911, _cvpt_1912, _cvpt_1913, _cvpt_1914, 
            _cvpt_1915, _cvpt_1916, _cvpt_1917, _cvpt_1918, _cvpt_1919, 
            _cvpt_1920, _cvpt_1921, _cvpt_1922, _cvpt_1923, _cvpt_1924, 
            _cvpt_1925, _cvpt_1926, _cvpt_1927, _cvpt_1928, _cvpt_1929, 
            _cvpt_1930, _cvpt_1931, _cvpt_1932, _cvpt_1933, _cvpt_1934, 
            _cvpt_1935, _cvpt_1936, _cvpt_1937, _cvpt_1938, _cvpt_1939, 
            _cvpt_1940, _cvpt_1941, _cvpt_1942, _cvpt_1943, _cvpt_1944, 
            _cvpt_1945, _cvpt_1946, _cvpt_1947, _cvpt_1948, _cvpt_1949, 
            _cvpt_1950, _cvpt_1951, _cvpt_1952, _cvpt_1953, _cvpt_1954, 
            _cvpt_1955, _cvpt_1956, _cvpt_1957, _cvpt_1958, _cvpt_1959, 
            _cvpt_1960, _cvpt_1961, _cvpt_1962, _cvpt_1963, _cvpt_1964, 
            _cvpt_1965, _cvpt_1966, _cvpt_1967, _cvpt_1968, _cvpt_1969, 
            _cvpt_1970, _cvpt_1971, _cvpt_1972, _cvpt_1973, _cvpt_1974, 
            _cvpt_1975, _cvpt_1976, _cvpt_1977, _cvpt_1978, _cvpt_1979, 
            _cvpt_1980, _cvpt_1981, _cvpt_1982, _cvpt_1983, _cvpt_1984, 
            _cvpt_1985, _cvpt_1986, _cvpt_1987, _cvpt_1988, _cvpt_1989, 
            _cvpt_1990, _cvpt_1991, _cvpt_1992, _cvpt_1993, _cvpt_1994, 
            _cvpt_1995, _cvpt_1996, _cvpt_1997, _cvpt_1998, _cvpt_1999, 
            _cvpt_2000, _cvpt_2001, _cvpt_2002, _cvpt_2003, _cvpt_2004, 
            _cvpt_2005, _cvpt_2006, _cvpt_2007, _cvpt_2008, _cvpt_2009, 
            _cvpt_2010, _cvpt_2011, _cvpt_2012, _cvpt_2013, _cvpt_2014, 
            _cvpt_2015, _cvpt_2016, _cvpt_2017, _cvpt_2018, _cvpt_2019, 
            _cvpt_2020, _cvpt_2021, _cvpt_2022, _cvpt_2023, _cvpt_2024, 
            _cvpt_2025, _cvpt_2026, _cvpt_2027, _cvpt_2028, _cvpt_2029, 
            _cvpt_2030, _cvpt_2031, _cvpt_2032, _cvpt_2033, _cvpt_2034, 
            _cvpt_2035, _cvpt_2036, _cvpt_2037, _cvpt_2038, _cvpt_2039, 
            _cvpt_2040, _cvpt_2041, _cvpt_2042, _cvpt_2043, _cvpt_2044, 
            _cvpt_2045, _cvpt_2046, _cvpt_2047, _cvpt_2048, _cvpt_2049, 
            _cvpt_2050, _cvpt_2051, _cvpt_2052, _cvpt_2053, _cvpt_2054, 
            _cvpt_2055, _cvpt_2056, _cvpt_2057, _cvpt_2058, _cvpt_2059, 
            _cvpt_2060, _cvpt_2061, _cvpt_2062, _cvpt_2063, _cvpt_2064, 
            _cvpt_2065, _cvpt_2066, _cvpt_2067, _cvpt_2068, _cvpt_2069, 
            _cvpt_2070, _cvpt_2071, _cvpt_2072, _cvpt_2073, _cvpt_2074, 
            _cvpt_2075, _cvpt_2076, _cvpt_2077, _cvpt_2078, _cvpt_2079, 
            _cvpt_2080, _cvpt_2081, _cvpt_2082, _cvpt_2083, _cvpt_2084, 
            _cvpt_2085, _cvpt_2086, _cvpt_2087, _cvpt_2088, _cvpt_2089, 
            _cvpt_2090, _cvpt_2091, _cvpt_2092, _cvpt_2093, _cvpt_2094, 
            _cvpt_2095, _cvpt_2096, _cvpt_2097, _cvpt_2098, _cvpt_2099, 
            _cvpt_2100, _cvpt_2101, _cvpt_2102, _cvpt_2103, _cvpt_2104, 
            _cvpt_2105, _cvpt_2106, _cvpt_2107, _cvpt_2108, _cvpt_2109, 
            _cvpt_2110, _cvpt_2111, _cvpt_2112, _cvpt_2113, _cvpt_2114, 
            _cvpt_2115, _cvpt_2116, _cvpt_2117, _cvpt_2118, _cvpt_2119, 
            _cvpt_2120, _cvpt_2121, _cvpt_2122, _cvpt_2123, _cvpt_2124, 
            _cvpt_2125, _cvpt_2126, _cvpt_2127, _cvpt_2128, _cvpt_2129, 
            _cvpt_2130, _cvpt_2131, _cvpt_2132, _cvpt_2133, _cvpt_2134, 
            _cvpt_2135, _cvpt_2136, _cvpt_2137, _cvpt_2138, _cvpt_2139, 
            _cvpt_2140, _cvpt_2141, _cvpt_2142, _cvpt_2143, _cvpt_2144, 
            _cvpt_2145, _cvpt_2146, _cvpt_2147, _cvpt_2148, _cvpt_2149, 
            _cvpt_2150, _cvpt_2151, _cvpt_2152, _cvpt_2153, _cvpt_2154, 
            _cvpt_2155, _cvpt_2156, _cvpt_2157, _cvpt_2158, _cvpt_2159, 
            _cvpt_2160, _cvpt_2161, _cvpt_2162, _cvpt_2163, _cvpt_2164, 
            _cvpt_2165, _cvpt_2166, _cvpt_2167, _cvpt_2168, _cvpt_2169, 
            _cvpt_2170, _cvpt_2171, _cvpt_2172, _cvpt_2173, _cvpt_2174, 
            _cvpt_2175, _cvpt_2176, _cvpt_2177, _cvpt_2178, _cvpt_2179, 
            _cvpt_2180, _cvpt_2181, _cvpt_2182, _cvpt_2183, _cvpt_2184, 
            _cvpt_2185, _cvpt_2186, _cvpt_2187, _cvpt_2188, _cvpt_2189, 
            _cvpt_2190, _cvpt_2191, _cvpt_2192, _cvpt_2193, _cvpt_2194, 
            _cvpt_2195, _cvpt_2196, _cvpt_2197, _cvpt_2198, _cvpt_2199, 
            _cvpt_2200, _cvpt_2201, _cvpt_2202, _cvpt_2203, _cvpt_2204, 
            _cvpt_2205, _cvpt_2206, _cvpt_2207, _cvpt_2208, _cvpt_2209, 
            _cvpt_2210, _cvpt_2211, _cvpt_2212, _cvpt_2213, _cvpt_2214, 
            _cvpt_2215, _cvpt_2216, _cvpt_2217, _cvpt_2218, _cvpt_2219, 
            _cvpt_2220, _cvpt_2221, _cvpt_2222, _cvpt_2223, _cvpt_2224, 
            _cvpt_2225, _cvpt_2226, _cvpt_2227, _cvpt_2228, _cvpt_2229, 
            _cvpt_2230, _cvpt_2231, _cvpt_2232, _cvpt_2233, _cvpt_2234, 
            _cvpt_2235, _cvpt_2236, _cvpt_2237, _cvpt_2238, _cvpt_2239, 
            _cvpt_2240, _cvpt_2241, _cvpt_2242, _cvpt_2243, _cvpt_2244, 
            _cvpt_2245, _cvpt_2246, _cvpt_2247, _cvpt_2248, _cvpt_2249, 
            _cvpt_2250, _cvpt_2251, _cvpt_2252, _cvpt_2253, _cvpt_2254, 
            _cvpt_2255, _cvpt_2256, _cvpt_2257, _cvpt_2258, _cvpt_2259, 
            _cvpt_2260, _cvpt_2261, _cvpt_2262, _cvpt_2263, _cvpt_2264, 
            _cvpt_2265, _cvpt_2266, _cvpt_2267, _cvpt_2268, _cvpt_2269, 
            _cvpt_2270, _cvpt_2271, _cvpt_2272, _cvpt_2273, _cvpt_2274, 
            _cvpt_2275, _cvpt_2276, _cvpt_2277, _cvpt_2278, _cvpt_2279, 
            _cvpt_2280, _cvpt_2281, _cvpt_2282, _cvpt_2283, _cvpt_2284, 
            _cvpt_2285, _cvpt_2286, _cvpt_2287, _cvpt_2288, _cvpt_2289, 
            _cvpt_2290, _cvpt_2291, _cvpt_2292, _cvpt_2293, _cvpt_2294, 
            _cvpt_2295, _cvpt_2296, _cvpt_2297, _cvpt_2298, _cvpt_2299, 
            _cvpt_2300, _cvpt_2301, _cvpt_2302, _cvpt_2303, _cvpt_2304, 
            _cvpt_2305, _cvpt_2306, _cvpt_2307, _cvpt_2308, _cvpt_2309, 
            _cvpt_2310, _cvpt_2311, _cvpt_2312, _cvpt_2313, _cvpt_2314, 
            _cvpt_2315, _cvpt_2316, _cvpt_2317, _cvpt_2318, _cvpt_2319, 
            _cvpt_2320, _cvpt_2321, _cvpt_2322, _cvpt_2323, _cvpt_2324, 
            _cvpt_2325, _cvpt_2326, _cvpt_2327, _cvpt_2328, _cvpt_2329, 
            _cvpt_2330, _cvpt_2331, _cvpt_2332, _cvpt_2333, _cvpt_2334, 
            _cvpt_2335, _cvpt_2336, _cvpt_2337, _cvpt_2338, _cvpt_2339, 
            _cvpt_2340, _cvpt_2341, _cvpt_2342, _cvpt_2343, _cvpt_2344, 
            _cvpt_2345, _cvpt_2346, _cvpt_2347, _cvpt_2348, _cvpt_2349, 
            _cvpt_2350, _cvpt_2351, _cvpt_2352, _cvpt_2353, _cvpt_2354, 
            _cvpt_2355, _cvpt_2356, _cvpt_2357, _cvpt_2358, _cvpt_2359, 
            _cvpt_2360, _cvpt_2361, _cvpt_2362, _cvpt_2363, _cvpt_2364, 
            _cvpt_2365, _cvpt_2366, _cvpt_2367, _cvpt_2368, _cvpt_2369, 
            _cvpt_2370, _cvpt_2371, _cvpt_2372, _cvpt_2373, _cvpt_2374, 
            _cvpt_2375, _cvpt_2376, _cvpt_2377, _cvpt_2378, _cvpt_2379, 
            _cvpt_2380, _cvpt_2381, _cvpt_2382, _cvpt_2383, _cvpt_2384, 
            _cvpt_2385, _cvpt_2386, _cvpt_2387, _cvpt_2388, _cvpt_2389, 
            _cvpt_2390, _cvpt_2391, _cvpt_2392, _cvpt_2393, _cvpt_2394, 
            _cvpt_2395, _cvpt_2396, _cvpt_2397, _cvpt_2398, _cvpt_2399, 
            _cvpt_2400, _cvpt_2401, _cvpt_2402, _cvpt_2403, _cvpt_2404, 
            _cvpt_2405, _cvpt_2406, _cvpt_2407, _cvpt_2408, _cvpt_2409, 
            _cvpt_2410, _cvpt_2411, _cvpt_2412, _cvpt_2413, _cvpt_2414, 
            _cvpt_2415, _cvpt_2416, _cvpt_2417, _cvpt_2418, _cvpt_2419, 
            _cvpt_2420, _cvpt_2421, _cvpt_2422, _cvpt_2423, _cvpt_2424, 
            _cvpt_2425, _cvpt_2426, _cvpt_2427, _cvpt_2428, _cvpt_2429, 
            _cvpt_2430, _cvpt_2431, _cvpt_2432, _cvpt_2433, _cvpt_2434, 
            _cvpt_2435, _cvpt_2436, _cvpt_2437, _cvpt_2438, _cvpt_2439, 
            _cvpt_2440, _cvpt_2441, _cvpt_2442, _cvpt_2443, _cvpt_2444, 
            _cvpt_2445, _cvpt_2446, _cvpt_2447, _cvpt_2448, _cvpt_2449, 
            _cvpt_2450, _cvpt_2451, _cvpt_2452, _cvpt_2453, _cvpt_2454, 
            _cvpt_2455, _cvpt_2456, _cvpt_2457, _cvpt_2458, _cvpt_2459, 
            _cvpt_2460, _cvpt_2461, _cvpt_2462, _cvpt_2463, _cvpt_2464, 
            _cvpt_2465, _cvpt_2466, _cvpt_2467, _cvpt_2468, _cvpt_2469, 
            _cvpt_2470, _cvpt_2471, _cvpt_2472, _cvpt_2473, _cvpt_2474, 
            _cvpt_2475, _cvpt_2476, _cvpt_2477, _cvpt_2478, _cvpt_2479, 
            _cvpt_2480, _cvpt_2481, _cvpt_2482, _cvpt_2483, _cvpt_2484, 
            _cvpt_2485, _cvpt_2486, _cvpt_2487, _cvpt_2488, _cvpt_2489, 
            _cvpt_2490, _cvpt_2491, _cvpt_2492, _cvpt_2493, _cvpt_2494, 
            _cvpt_2495, _cvpt_2496, _cvpt_2497, _cvpt_2498, _cvpt_2499, 
            _cvpt_2500, _cvpt_2501, _cvpt_2502, _cvpt_2503, _cvpt_2504, 
            _cvpt_2505, _cvpt_2506, _cvpt_2507, _cvpt_2508, _cvpt_2509, 
            _cvpt_2510, _cvpt_2511, _cvpt_2512, _cvpt_2513, _cvpt_2514, 
            _cvpt_2515, _cvpt_2516, _cvpt_2517, _cvpt_2518, _cvpt_2519, 
            _cvpt_2520, _cvpt_2521, _cvpt_2522, _cvpt_2523, _cvpt_2524, 
            _cvpt_2525, _cvpt_2526, _cvpt_2527, _cvpt_2528, _cvpt_2529, 
            _cvpt_2530, _cvpt_2531, _cvpt_2532, _cvpt_2533, _cvpt_2534, 
            _cvpt_2535, _cvpt_2536, _cvpt_2537, _cvpt_2538, _cvpt_2539, 
            _cvpt_2540, _cvpt_2541, _cvpt_2542, _cvpt_2543, _cvpt_2544, 
            _cvpt_2545, _cvpt_2546, _cvpt_2547, _cvpt_2548, _cvpt_2549, 
            _cvpt_2550, _cvpt_2551, _cvpt_2552, _cvpt_2553, _cvpt_2554, 
            _cvpt_2555, _cvpt_2556, _cvpt_2557, _cvpt_2558, _cvpt_2559, 
            _cvpt_2560, _cvpt_2561, _cvpt_2562, _cvpt_2563, _cvpt_2564, 
            _cvpt_2565, _cvpt_2566, _cvpt_2567, _cvpt_2568, _cvpt_2569, 
            _cvpt_2570, _cvpt_2571, _cvpt_2572, _cvpt_2573, _cvpt_2574, 
            _cvpt_2575, _cvpt_2576, _cvpt_2577, _cvpt_2578, _cvpt_2579, 
            _cvpt_2580, _cvpt_2581, _cvpt_2582, _cvpt_2583, _cvpt_2584, 
            _cvpt_2585, _cvpt_2586, _cvpt_2587, _cvpt_2588, _cvpt_2589, 
            _cvpt_2590, _cvpt_2591, _cvpt_2592, _cvpt_2593, _cvpt_2594, 
            _cvpt_2595, _cvpt_2596, _cvpt_2597, _cvpt_2598, _cvpt_2599, 
            _cvpt_2600, _cvpt_2601, _cvpt_2602, _cvpt_2603, _cvpt_2604, 
            _cvpt_2605, _cvpt_2606, _cvpt_2607, _cvpt_2608, _cvpt_2609, 
            _cvpt_2610, _cvpt_2611, _cvpt_2612, _cvpt_2613, _cvpt_2614, 
            _cvpt_2615, _cvpt_2616, _cvpt_2617, _cvpt_2618, _cvpt_2619, 
            _cvpt_2620, _cvpt_2621, _cvpt_2622, _cvpt_2623, _cvpt_2624, 
            _cvpt_2625, _cvpt_2626, _cvpt_2627, _cvpt_2628, _cvpt_2629, 
            _cvpt_2630, _cvpt_2631, _cvpt_2632, _cvpt_2633, _cvpt_2634, 
            _cvpt_2635, _cvpt_2636, _cvpt_2637, _cvpt_2638, _cvpt_2639, 
            _cvpt_2640, _cvpt_2641, _cvpt_2642, _cvpt_2643, _cvpt_2644, 
            _cvpt_2645, _cvpt_2646, _cvpt_2647, _cvpt_2648, _cvpt_2649, 
            _cvpt_2650, _cvpt_2651, _cvpt_2652, _cvpt_2653, _cvpt_2654, 
            _cvpt_2655, _cvpt_2656, _cvpt_2657, _cvpt_2658, _cvpt_2659, 
            _cvpt_2660, _cvpt_2661, _cvpt_2662, _cvpt_2663, _cvpt_2664, 
            _cvpt_2665, _cvpt_2666, _cvpt_2667, _cvpt_2668, _cvpt_2669, 
            _cvpt_2670, _cvpt_2671, _cvpt_2672, _cvpt_2673, _cvpt_2674, 
            _cvpt_2675, _cvpt_2676, _cvpt_2677, _cvpt_2678, _cvpt_2679, 
            _cvpt_2680, _cvpt_2681, _cvpt_2682, _cvpt_2683, _cvpt_2684, 
            _cvpt_2685, _cvpt_2686, _cvpt_2687, _cvpt_2688, _cvpt_2689, 
            _cvpt_2690, _cvpt_2691, _cvpt_2692, _cvpt_2693, _cvpt_2694, 
            _cvpt_2695, _cvpt_2696, _cvpt_2697, _cvpt_2698, _cvpt_2699, 
            _cvpt_2700, _cvpt_2701, _cvpt_2702, _cvpt_2703, _cvpt_2704, 
            _cvpt_2705, _cvpt_2706, _cvpt_2707, _cvpt_2708, _cvpt_2709, 
            _cvpt_2710, _cvpt_2711, _cvpt_2712, _cvpt_2713, _cvpt_2714, 
            _cvpt_2715, _cvpt_2716, _cvpt_2717, _cvpt_2718, _cvpt_2719, 
            _cvpt_2720, _cvpt_2721, _cvpt_2722, _cvpt_2723, _cvpt_2724, 
            _cvpt_2725, _cvpt_2726, _cvpt_2727, _cvpt_2728, _cvpt_2729, 
            _cvpt_2730, _cvpt_2731, _cvpt_2732, _cvpt_2733, _cvpt_2734, 
            _cvpt_2735, _cvpt_2736, _cvpt_2737, _cvpt_2738, _cvpt_2739, 
            _cvpt_2740, _cvpt_2741, _cvpt_2742, _cvpt_2743, _cvpt_2744, 
            _cvpt_2745, _cvpt_2746, _cvpt_2747, _cvpt_2748, _cvpt_2749, 
            _cvpt_2750, _cvpt_2751, _cvpt_2752, _cvpt_2753, _cvpt_2754, 
            _cvpt_2755, _cvpt_2756, _cvpt_2757, _cvpt_2758, _cvpt_2759, 
            _cvpt_2760, _cvpt_2761, _cvpt_2762, _cvpt_2763, _cvpt_2764, 
            _cvpt_2765, _cvpt_2766, _cvpt_2767, _cvpt_2768, _cvpt_2769, 
            _cvpt_2770, _cvpt_2771, _cvpt_2772, _cvpt_2773, _cvpt_2774, 
            _cvpt_2775, _cvpt_2776, _cvpt_2777, _cvpt_2778, _cvpt_2779, 
            _cvpt_2780, _cvpt_2781, _cvpt_2782, _cvpt_2783, _cvpt_2784, 
            _cvpt_2785, _cvpt_2786, _cvpt_2787, _cvpt_2788, _cvpt_2789, 
            _cvpt_2790, _cvpt_2791, _cvpt_2792, _cvpt_2793, _cvpt_2794, 
            _cvpt_2795, _cvpt_2796, _cvpt_2797, _cvpt_2798, _cvpt_2799, 
            _cvpt_2800, _cvpt_2801, _cvpt_2802, _cvpt_2803, _cvpt_2804, 
            _cvpt_2805, _cvpt_2806, _cvpt_2807, _cvpt_2808, _cvpt_2809, 
            _cvpt_2810, _cvpt_2811, _cvpt_2812, _cvpt_2813, _cvpt_2814, 
            _cvpt_2815, _cvpt_2816, _cvpt_2817, _cvpt_2818, _cvpt_2819, 
            _cvpt_2820, _cvpt_2821, _cvpt_2822, _cvpt_2823, _cvpt_2824, 
            _cvpt_2825, _cvpt_2826, _cvpt_2827, _cvpt_2828, _cvpt_2829, 
            _cvpt_2830, _cvpt_2831, _cvpt_2832, _cvpt_2833, _cvpt_2834, 
            _cvpt_2835, _cvpt_2836, _cvpt_2837, _cvpt_2838, _cvpt_2839, 
            _cvpt_2840, _cvpt_2841, _cvpt_2842, _cvpt_2843, _cvpt_2844, 
            _cvpt_2845, _cvpt_2846, _cvpt_2847, _cvpt_2848, _cvpt_2849, 
            _cvpt_2850, _cvpt_2851, _cvpt_2852, _cvpt_2853, _cvpt_2854, 
            _cvpt_2855, _cvpt_2856, _cvpt_2857, _cvpt_2858, _cvpt_2859, 
            _cvpt_2860, _cvpt_2861, _cvpt_2862, _cvpt_2863, _cvpt_2864, 
            _cvpt_2865, _cvpt_2866, _cvpt_2867, _cvpt_2868, _cvpt_2869, 
            _cvpt_2870, _cvpt_2871, _cvpt_2872, _cvpt_2873, _cvpt_2874, 
            _cvpt_2875, _cvpt_2876, _cvpt_2877, _cvpt_2878, _cvpt_2879, 
            _cvpt_2880, _cvpt_2881, _cvpt_2882, _cvpt_2883, _cvpt_2884, 
            _cvpt_2885, _cvpt_2886, _cvpt_2887, _cvpt_2888, _cvpt_2889, 
            _cvpt_2890, _cvpt_2891, _cvpt_2892, _cvpt_2893, _cvpt_2894, 
            _cvpt_2895, _cvpt_2896, _cvpt_2897, _cvpt_2898, _cvpt_2899, 
            _cvpt_2900, _cvpt_2901, _cvpt_2902, _cvpt_2903, _cvpt_2904, 
            _cvpt_2905, _cvpt_2906, _cvpt_2907, _cvpt_2908, _cvpt_2909, 
            _cvpt_2910, _cvpt_2911, _cvpt_2912, _cvpt_2913, _cvpt_2914, 
            _cvpt_2915, _cvpt_2916, _cvpt_2917, _cvpt_2918, _cvpt_2919, 
            _cvpt_2920, _cvpt_2921, _cvpt_2922, _cvpt_2923, _cvpt_2924, 
            _cvpt_2925, _cvpt_2926, _cvpt_2927, _cvpt_2928, _cvpt_2929, 
            _cvpt_2930, _cvpt_2931, _cvpt_2932, _cvpt_2933, _cvpt_2934, 
            _cvpt_2935, _cvpt_2936, _cvpt_2937, _cvpt_2938, _cvpt_2939, 
            _cvpt_2940, _cvpt_2941, _cvpt_2942, _cvpt_2943, _cvpt_2944, 
            _cvpt_2945, _cvpt_2946, _cvpt_2947, _cvpt_2948, _cvpt_2949, 
            _cvpt_2950, _cvpt_2951, _cvpt_2952, _cvpt_2953, _cvpt_2954, 
            _cvpt_2955, _cvpt_2956, _cvpt_2957, _cvpt_2958, _cvpt_2959, 
            _cvpt_2960, _cvpt_2961, _cvpt_2962, _cvpt_2963, _cvpt_2964, 
            _cvpt_2965, _cvpt_2966, _cvpt_2967, _cvpt_2968, _cvpt_2969, 
            _cvpt_2970, _cvpt_2971, _cvpt_2972, _cvpt_2973, _cvpt_2974, 
            _cvpt_2975, _cvpt_2976, _cvpt_2977, _cvpt_2978, _cvpt_2979, 
            _cvpt_2980, _cvpt_2981, _cvpt_2982, _cvpt_2983, _cvpt_2984, 
            _cvpt_2985, _cvpt_2986, _cvpt_2987, _cvpt_2988, _cvpt_2989, 
            _cvpt_2990, _cvpt_2991, _cvpt_2992, _cvpt_2993, _cvpt_2994, 
            _cvpt_2995, _cvpt_2996, _cvpt_2997, _cvpt_2998, _cvpt_2999, 
            _cvpt_3000, _cvpt_3001, _cvpt_3002, _cvpt_3003, _cvpt_3004, 
            _cvpt_3005, _cvpt_3006, _cvpt_3007, _cvpt_3008, _cvpt_3009, 
            _cvpt_3010, _cvpt_3011, _cvpt_3012, _cvpt_3013, _cvpt_3014, 
            _cvpt_3015, _cvpt_3016, _cvpt_3017, _cvpt_3018, _cvpt_3019, 
            _cvpt_3020, _cvpt_3021, _cvpt_3022, _cvpt_3023, _cvpt_3024, 
            _cvpt_3025, _cvpt_3026, _cvpt_3027, _cvpt_3028, _cvpt_3029, 
            _cvpt_3030, _cvpt_3031, _cvpt_3032, _cvpt_3033, _cvpt_3034, 
            _cvpt_3035, _cvpt_3036, _cvpt_3037, _cvpt_3038, _cvpt_3039, 
            _cvpt_3040, _cvpt_3041, _cvpt_3042, _cvpt_3043, _cvpt_3044, 
            _cvpt_3045, _cvpt_3046, _cvpt_3047, _cvpt_3048, _cvpt_3049, 
            _cvpt_3050, _cvpt_3051, _cvpt_3052, _cvpt_3053, _cvpt_3054, 
            _cvpt_3055, _cvpt_3056, _cvpt_3057, _cvpt_3058, _cvpt_3059, 
            _cvpt_3060, _cvpt_3061, _cvpt_3062, _cvpt_3063, _cvpt_3064, 
            _cvpt_3065, _cvpt_3066, _cvpt_3067, _cvpt_3068, _cvpt_3069, 
            _cvpt_3070, _cvpt_3071, _cvpt_3072, _cvpt_3073, _cvpt_3074, 
            _cvpt_3075, _cvpt_3076, _cvpt_3077, _cvpt_3078, _cvpt_3079, 
            _cvpt_3080, _cvpt_3081, _cvpt_3082, _cvpt_3083, _cvpt_3084, 
            _cvpt_3085, _cvpt_3086, _cvpt_3087, _cvpt_3088, _cvpt_3089, 
            _cvpt_3090, _cvpt_3091, _cvpt_3092, _cvpt_3093, _cvpt_3094, 
            _cvpt_3095, _cvpt_3096, _cvpt_3097, _cvpt_3098, _cvpt_3099, 
            _cvpt_3100, _cvpt_3101, _cvpt_3102, _cvpt_3103, _cvpt_3104, 
            _cvpt_3105, _cvpt_3106, _cvpt_3107, _cvpt_3108, _cvpt_3109, 
            _cvpt_3110, _cvpt_3111, _cvpt_3112, _cvpt_3113, _cvpt_3114, 
            _cvpt_3115, _cvpt_3116, _cvpt_3117, _cvpt_3118, _cvpt_3119, 
            _cvpt_3120, _cvpt_3121, _cvpt_3122, _cvpt_3123, _cvpt_3124, 
            _cvpt_3125, _cvpt_3126, _cvpt_3127, _cvpt_3128, _cvpt_3129, 
            _cvpt_3130, _cvpt_3131, _cvpt_3132, _cvpt_3133, _cvpt_3134, 
            _cvpt_3135, _cvpt_3136, _cvpt_3137, _cvpt_3138, _cvpt_3139, 
            _cvpt_3140, _cvpt_3141, _cvpt_3142, _cvpt_3143, _cvpt_3144, 
            _cvpt_3145, _cvpt_3146, _cvpt_3147, _cvpt_3148, _cvpt_3149, 
            _cvpt_3150, _cvpt_3151, _cvpt_3152, _cvpt_3153, _cvpt_3154, 
            _cvpt_3155, _cvpt_3156, _cvpt_3157, _cvpt_3158, _cvpt_3159, 
            _cvpt_3160, _cvpt_3161, _cvpt_3162, _cvpt_3163, _cvpt_3164, 
            _cvpt_3165, _cvpt_3166, _cvpt_3167, _cvpt_3168, _cvpt_3169, 
            _cvpt_3170, _cvpt_3171, _cvpt_3172, _cvpt_3173, _cvpt_3174, 
            _cvpt_3175, _cvpt_3176, _cvpt_3177, _cvpt_3178, _cvpt_3179, 
            _cvpt_3180, _cvpt_3181, _cvpt_3182, _cvpt_3183, _cvpt_3184, 
            _cvpt_3185, _cvpt_3186, _cvpt_3187, _cvpt_3188, _cvpt_3189, 
            _cvpt_3190, _cvpt_3191, _cvpt_3192, _cvpt_3193, _cvpt_3194, 
            _cvpt_3195, _cvpt_3196, _cvpt_3197, _cvpt_3198, _cvpt_3199, 
            _cvpt_3200, _cvpt_3201, _cvpt_3202, _cvpt_3203, _cvpt_3204, 
            _cvpt_3205, _cvpt_3206, _cvpt_3207, _cvpt_3208, _cvpt_3209, 
            _cvpt_3210, _cvpt_3211, _cvpt_3212, _cvpt_3213, _cvpt_3214, 
            _cvpt_3215, _cvpt_3216, _cvpt_3217, _cvpt_3218, _cvpt_3219, 
            _cvpt_3220, _cvpt_3221, _cvpt_3222, _cvpt_3223, _cvpt_3224, 
            _cvpt_3225, _cvpt_3226, _cvpt_3227, _cvpt_3228, _cvpt_3229, 
            _cvpt_3230, _cvpt_3231, _cvpt_3232, _cvpt_3233, _cvpt_3234, 
            _cvpt_3235, _cvpt_3236, _cvpt_3237, _cvpt_3238, _cvpt_3239, 
            _cvpt_3240, _cvpt_3241, _cvpt_3242, _cvpt_3243, _cvpt_3244, 
            _cvpt_3245, _cvpt_3246, _cvpt_3247, _cvpt_3248, _cvpt_3249, 
            _cvpt_3250, _cvpt_3251, _cvpt_3252, _cvpt_3253, _cvpt_3254, 
            _cvpt_3255, _cvpt_3256, _cvpt_3257, _cvpt_3258, _cvpt_3259, 
            _cvpt_3260, _cvpt_3261, _cvpt_3262, _cvpt_3263, _cvpt_3264, 
            _cvpt_3265, _cvpt_3266, _cvpt_3267, _cvpt_3268, _cvpt_3269, 
            _cvpt_3270, _cvpt_3271, _cvpt_3272, _cvpt_3273, _cvpt_3274, 
            _cvpt_3275, _cvpt_3276, _cvpt_3277, _cvpt_3278, _cvpt_3279, 
            _cvpt_3280, _cvpt_3281, _cvpt_3282, _cvpt_3283, _cvpt_3284, 
            _cvpt_3285, _cvpt_3286, _cvpt_3287, _cvpt_3288, _cvpt_3289, 
            _cvpt_3290, _cvpt_3291, _cvpt_3292, _cvpt_3293, _cvpt_3294, 
            _cvpt_3295, _cvpt_3296, _cvpt_3297, _cvpt_3298, _cvpt_3299, 
            _cvpt_3300, _cvpt_3301, _cvpt_3302, _cvpt_3303, _cvpt_3304, 
            _cvpt_3305, _cvpt_3306, _cvpt_3307, _cvpt_3308, _cvpt_3309, 
            _cvpt_3310, _cvpt_3311, _cvpt_3312, _cvpt_3313, _cvpt_3314, 
            _cvpt_3315, _cvpt_3316, _cvpt_3317, _cvpt_3318, _cvpt_3319, 
            _cvpt_3320, _cvpt_3321, _cvpt_3322, _cvpt_3323, _cvpt_3324, 
            _cvpt_3325, _cvpt_3326, _cvpt_3327, _cvpt_3328, _cvpt_3329, 
            _cvpt_3330, _cvpt_3331, _cvpt_3332, _cvpt_3333, _cvpt_3334, 
            _cvpt_3335, _cvpt_3336, _cvpt_3337, _cvpt_3338, _cvpt_3339, 
            _cvpt_3340, _cvpt_3341, _cvpt_3342, _cvpt_3343, _cvpt_3344, 
            _cvpt_3345, _cvpt_3346, _cvpt_3347, _cvpt_3348, _cvpt_3349, 
            _cvpt_3350, _cvpt_3351, _cvpt_3352, _cvpt_3353, _cvpt_3354, 
            _cvpt_3355, _cvpt_3356, _cvpt_3357, _cvpt_3358, _cvpt_3359, 
            _cvpt_3360, _cvpt_3361, _cvpt_3362, _cvpt_3363, _cvpt_3364, 
            _cvpt_3365, _cvpt_3366, _cvpt_3367, _cvpt_3368, _cvpt_3369, 
            _cvpt_3370, _cvpt_3371, _cvpt_3372, _cvpt_3373, _cvpt_3374, 
            _cvpt_3375, _cvpt_3376, _cvpt_3377, _cvpt_3378, _cvpt_3379, 
            _cvpt_3380, _cvpt_3381, _cvpt_3382, _cvpt_3383, _cvpt_3384, 
            _cvpt_3385, _cvpt_3386, _cvpt_3387, _cvpt_3388, _cvpt_3389, 
            _cvpt_3390, _cvpt_3391, _cvpt_3392, _cvpt_3393, _cvpt_3394, 
            _cvpt_3395, _cvpt_3396, _cvpt_3397, _cvpt_3398, _cvpt_3399, 
            _cvpt_3400, _cvpt_3401, _cvpt_3402, _cvpt_3403, _cvpt_3404, 
            _cvpt_3405, _cvpt_3406, _cvpt_3407, _cvpt_3408, _cvpt_3409, 
            _cvpt_3410, _cvpt_3411, _cvpt_3412, _cvpt_3413, _cvpt_3414, 
            _cvpt_3415, _cvpt_3416, _cvpt_3417, _cvpt_3418, _cvpt_3419, 
            _cvpt_3420, _cvpt_3421, _cvpt_3422, _cvpt_3423, _cvpt_3424, 
            _cvpt_3425, _cvpt_3426, _cvpt_3427, _cvpt_3428, _cvpt_3429, 
            _cvpt_3430, _cvpt_3431, _cvpt_3432, _cvpt_3433, _cvpt_3434, 
            _cvpt_3435, _cvpt_3436, _cvpt_3437, _cvpt_3438, _cvpt_3439, 
            _cvpt_3440, _cvpt_3441, _cvpt_3442, _cvpt_3443, _cvpt_3444, 
            _cvpt_3445, _cvpt_3446, _cvpt_3447, _cvpt_3448, _cvpt_3449, 
            _cvpt_3450, _cvpt_3451, _cvpt_3452, _cvpt_3453, _cvpt_3454, 
            _cvpt_3455, _cvpt_3456, _cvpt_3457, _cvpt_3458, _cvpt_3459, 
            _cvpt_3460, _cvpt_3461, _cvpt_3462, _cvpt_3463, _cvpt_3464, 
            _cvpt_3465, _cvpt_3466, _cvpt_3467, _cvpt_3468, _cvpt_3469, 
            _cvpt_3470, _cvpt_3471, _cvpt_3472, _cvpt_3473, _cvpt_3474, 
            _cvpt_3475, _cvpt_3476, _cvpt_3477, _cvpt_3478, _cvpt_3479, 
            _cvpt_3480, _cvpt_3481, _cvpt_3482, _cvpt_3483, _cvpt_3484, 
            _cvpt_3485, _cvpt_3486, _cvpt_3487, _cvpt_3488, _cvpt_3489, 
            _cvpt_3490, _cvpt_3491, _cvpt_3492, _cvpt_3493, _cvpt_3494, 
            _cvpt_3495, _cvpt_3496, _cvpt_3497, _cvpt_3498, _cvpt_3499, 
            _cvpt_3500, _cvpt_3501, _cvpt_3502, _cvpt_3503, _cvpt_3504, 
            _cvpt_3505, _cvpt_3506, _cvpt_3507, _cvpt_3508, _cvpt_3509, 
            _cvpt_3510, _cvpt_3511, _cvpt_3512, _cvpt_3513, _cvpt_3514, 
            _cvpt_3515, _cvpt_3516, _cvpt_3517, _cvpt_3518, _cvpt_3519, 
            _cvpt_3520, _cvpt_3521, _cvpt_3522, _cvpt_3523, _cvpt_3524, 
            _cvpt_3525, _cvpt_3526, _cvpt_3527, _cvpt_3528, _cvpt_3529, 
            _cvpt_3530, _cvpt_3531, _cvpt_3532, _cvpt_3533, _cvpt_3534, 
            _cvpt_3535, _cvpt_3536, _cvpt_3537, _cvpt_3538, _cvpt_3539, 
            _cvpt_3540, _cvpt_3541, _cvpt_3542, _cvpt_3543, _cvpt_3544, 
            _cvpt_3545, _cvpt_3546, _cvpt_3547, _cvpt_3548, _cvpt_3549, 
            _cvpt_3550, _cvpt_3551, _cvpt_3552, _cvpt_3553, _cvpt_3554, 
            _cvpt_3555, _cvpt_3556, _cvpt_3557, _cvpt_3558, _cvpt_3559, 
            _cvpt_3560, _cvpt_3561, _cvpt_3562, _cvpt_3563, _cvpt_3564, 
            _cvpt_3565, _cvpt_3566, _cvpt_3567, _cvpt_3568, _cvpt_3569, 
            _cvpt_3570, _cvpt_3571, _cvpt_3572, _cvpt_3573, _cvpt_3574, 
            _cvpt_3575, _cvpt_3576, _cvpt_3577, _cvpt_3578, _cvpt_3579, 
            _cvpt_3580, _cvpt_3581, _cvpt_3582, _cvpt_3583, _cvpt_3584, 
            _cvpt_3585, _cvpt_3586, _cvpt_3587, _cvpt_3588, _cvpt_3589, 
            _cvpt_3590, _cvpt_3591, _cvpt_3592, _cvpt_3593, _cvpt_3594, 
            _cvpt_3595, _cvpt_3596, _cvpt_3597, _cvpt_3598, _cvpt_3599, 
            _cvpt_3600, _cvpt_3601, _cvpt_3602, _cvpt_3603, _cvpt_3604, 
            _cvpt_3605, _cvpt_3606, _cvpt_3607, _cvpt_3608, _cvpt_3609, 
            _cvpt_3610, _cvpt_3611, _cvpt_3612, _cvpt_3613, _cvpt_3614, 
            _cvpt_3615, _cvpt_3616, _cvpt_3617, _cvpt_3618, _cvpt_3619, 
            _cvpt_3620, _cvpt_3621, _cvpt_3622, _cvpt_3623, _cvpt_3624, 
            _cvpt_3625, _cvpt_3626, _cvpt_3627, _cvpt_3628, _cvpt_3629, 
            _cvpt_3630, _cvpt_3631, _cvpt_3632, _cvpt_3633, _cvpt_3634, 
            _cvpt_3635, _cvpt_3636, _cvpt_3637, _cvpt_3638, _cvpt_3639, 
            _cvpt_3640, _cvpt_3641, _cvpt_3642, _cvpt_3643, _cvpt_3644, 
            _cvpt_3645, _cvpt_3646, _cvpt_3647, _cvpt_3648, _cvpt_3649, 
            _cvpt_3650, _cvpt_3651, _cvpt_3652, _cvpt_3653, _cvpt_3654, 
            _cvpt_3655, _cvpt_3656, _cvpt_3657, _cvpt_3658, _cvpt_3659, 
            _cvpt_3660, _cvpt_3661, _cvpt_3662, _cvpt_3663, _cvpt_3664, 
            _cvpt_3665, _cvpt_3666, _cvpt_3667, _cvpt_3668, _cvpt_3669, 
            _cvpt_3670, _cvpt_3671, _cvpt_3672, _cvpt_3673, _cvpt_3674, 
            _cvpt_3675, _cvpt_3676, _cvpt_3677, _cvpt_3678, _cvpt_3679, 
            _cvpt_3680, _cvpt_3681, _cvpt_3682, _cvpt_3683, _cvpt_3684, 
            _cvpt_3685, _cvpt_3686, _cvpt_3687, _cvpt_3688, _cvpt_3689, 
            _cvpt_3690, _cvpt_3691, _cvpt_3692, _cvpt_3693, _cvpt_3694, 
            _cvpt_3695, _cvpt_3696, _cvpt_3697, _cvpt_3698, _cvpt_3699, 
            _cvpt_3700, _cvpt_3701, _cvpt_3702, _cvpt_3703, _cvpt_3704, 
            _cvpt_3705, _cvpt_3706, _cvpt_3707, _cvpt_3708, _cvpt_3709, 
            _cvpt_3710, _cvpt_3711, _cvpt_3712, _cvpt_3713, _cvpt_3714, 
            _cvpt_3715, _cvpt_3716, _cvpt_3717, _cvpt_3718, _cvpt_3719, 
            _cvpt_3720, _cvpt_3721, _cvpt_3722, _cvpt_3723, _cvpt_3724, 
            _cvpt_3725, _cvpt_3726, _cvpt_3727, _cvpt_3728, _cvpt_3729, 
            _cvpt_3730, _cvpt_3731, _cvpt_3732, _cvpt_3733, _cvpt_3734, 
            _cvpt_3735, _cvpt_3736, _cvpt_3737, _cvpt_3738, _cvpt_3739, 
            _cvpt_3740, _cvpt_3741, _cvpt_3742, _cvpt_3743, _cvpt_3744, 
            _cvpt_3745, _cvpt_3746, _cvpt_3747, _cvpt_3748, _cvpt_3749, 
            _cvpt_3750, _cvpt_3751, _cvpt_3752, _cvpt_3753, _cvpt_3754, 
            _cvpt_3755, _cvpt_3756, _cvpt_3757, _cvpt_3758, _cvpt_3759, 
            _cvpt_3760, _cvpt_3761, _cvpt_3762, _cvpt_3763, _cvpt_3764, 
            _cvpt_3765, _cvpt_3766, _cvpt_3767, _cvpt_3768, _cvpt_3769, 
            _cvpt_3770, _cvpt_3771, _cvpt_3772, _cvpt_3773, _cvpt_3774, 
            _cvpt_3775, _cvpt_3776, _cvpt_3777, _cvpt_3778, _cvpt_3779, 
            _cvpt_3780, _cvpt_3781, _cvpt_3782, _cvpt_3783, _cvpt_3784, 
            _cvpt_3785, _cvpt_3786, _cvpt_3787, _cvpt_3788, _cvpt_3789, 
            _cvpt_3790, _cvpt_3791, _cvpt_3792, _cvpt_3793, _cvpt_3794, 
            _cvpt_3795, _cvpt_3796, _cvpt_3797, _cvpt_3798, _cvpt_3799, 
            _cvpt_3800, _cvpt_3801, _cvpt_3802, _cvpt_3803, _cvpt_3804, 
            _cvpt_3805, _cvpt_3806, _cvpt_3807, _cvpt_3808, _cvpt_3809, 
            _cvpt_3810, _cvpt_3811, _cvpt_3812, _cvpt_3813, _cvpt_3814, 
            _cvpt_3815, _cvpt_3816, _cvpt_3817, _cvpt_3818, _cvpt_3819, 
            _cvpt_3820, _cvpt_3821, _cvpt_3822, _cvpt_3823, _cvpt_3824, 
            _cvpt_3825, _cvpt_3826, _cvpt_3827, _cvpt_3828, _cvpt_3829, 
            _cvpt_3830, _cvpt_3831, _cvpt_3832, _cvpt_3833, _cvpt_3834, 
            _cvpt_3835, _cvpt_3836, _cvpt_3837, _cvpt_3838, _cvpt_3839, 
            _cvpt_3840, _cvpt_3841, _cvpt_3842, _cvpt_3843, _cvpt_3844, 
            _cvpt_3845, _cvpt_3846, _cvpt_3847, _cvpt_3848, _cvpt_3849, 
            _cvpt_3850, _cvpt_3851, _cvpt_3852, _cvpt_3853, _cvpt_3854, 
            _cvpt_3855, _cvpt_3856, _cvpt_3857, _cvpt_3858, _cvpt_3859, 
            _cvpt_3860, _cvpt_3861, _cvpt_3862, _cvpt_3863, _cvpt_3864, 
            _cvpt_3865, _cvpt_3866, _cvpt_3867, _cvpt_3868, _cvpt_3869, 
            _cvpt_3870, _cvpt_3871, _cvpt_3872, _cvpt_3873, _cvpt_3874, 
            _cvpt_3875, _cvpt_3876, _cvpt_3877, _cvpt_3878, _cvpt_3879, 
            _cvpt_3880, _cvpt_3881, _cvpt_3882, _cvpt_3883, _cvpt_3884, 
            _cvpt_3885, _cvpt_3886, _cvpt_3887, _cvpt_3888, _cvpt_3889, 
            _cvpt_3890, _cvpt_3891, _cvpt_3892, _cvpt_3893, _cvpt_3894, 
            _cvpt_3895, _cvpt_3896, _cvpt_3897, _cvpt_3898, _cvpt_3899, 
            _cvpt_3900, _cvpt_3901, _cvpt_3902, _cvpt_3903, _cvpt_3904, 
            _cvpt_3905, _cvpt_3906, _cvpt_3907, _cvpt_3908, _cvpt_3909, 
            _cvpt_3910, _cvpt_3911, _cvpt_3912, _cvpt_3913, _cvpt_3914, 
            _cvpt_3915, _cvpt_3916, _cvpt_3917, _cvpt_3918, _cvpt_3919, 
            _cvpt_3920, _cvpt_3921, _cvpt_3922, _cvpt_3923, _cvpt_3924, 
            _cvpt_3925, _cvpt_3926, _cvpt_3927, _cvpt_3928, _cvpt_3929, 
            _cvpt_3930, _cvpt_3931, _cvpt_3932, _cvpt_3933, _cvpt_3934, 
            _cvpt_3935, _cvpt_3936, _cvpt_3937, _cvpt_3938, _cvpt_3939, 
            _cvpt_3940, _cvpt_3941, _cvpt_3942, _cvpt_3943, _cvpt_3944, 
            _cvpt_3945, _cvpt_3946, _cvpt_3947, _cvpt_3948, _cvpt_3949, 
            _cvpt_3950, _cvpt_3951, _cvpt_3952, _cvpt_3953, _cvpt_3954, 
            _cvpt_3955, _cvpt_3956, _cvpt_3957, _cvpt_3958, _cvpt_3959, 
            _cvpt_3960, _cvpt_3961, _cvpt_3962, _cvpt_3963, _cvpt_3964, 
            _cvpt_3965, _cvpt_3966, _cvpt_3967, _cvpt_3968, _cvpt_3969, 
            _cvpt_3970, _cvpt_3971, _cvpt_3972, _cvpt_3973, _cvpt_3974, 
            _cvpt_3975, _cvpt_3976, _cvpt_3977, _cvpt_3978, _cvpt_3979, 
            _cvpt_3980, _cvpt_3981, _cvpt_3982, _cvpt_3983, _cvpt_3984, 
            _cvpt_3985, _cvpt_3986, _cvpt_3987, _cvpt_3988, _cvpt_3989, 
            _cvpt_3990, _cvpt_3991, _cvpt_3992, _cvpt_3993, _cvpt_3994, 
            _cvpt_3995, _cvpt_3996, _cvpt_3997, _cvpt_3998, _cvpt_3999, 
            _cvpt_4000, _cvpt_4001, _cvpt_4002, _cvpt_4003, _cvpt_4004, 
            _cvpt_4005, _cvpt_4006, _cvpt_4007, _cvpt_4008, _cvpt_4009, 
            _cvpt_4010, _cvpt_4011, _cvpt_4012, _cvpt_4013, _cvpt_4014, 
            _cvpt_4015, _cvpt_4016, _cvpt_4017, _cvpt_4018, _cvpt_4019, 
            _cvpt_4020, _cvpt_4021, _cvpt_4022, _cvpt_4023, _cvpt_4024, 
            _cvpt_4025, _cvpt_4026, _cvpt_4027, _cvpt_4028, _cvpt_4029, 
            _cvpt_4030, _cvpt_4031, _cvpt_4032, _cvpt_4033, _cvpt_4034, 
            _cvpt_4035, _cvpt_4036, _cvpt_4037, _cvpt_4038, _cvpt_4039, 
            _cvpt_4040, _cvpt_4041, _cvpt_4042, _cvpt_4043, _cvpt_4044, 
            _cvpt_4045, _cvpt_4046, _cvpt_4047, _cvpt_4048, _cvpt_4049, 
            _cvpt_4050, _cvpt_4051, _cvpt_4052, _cvpt_4053, _cvpt_4054, 
            _cvpt_4055, _cvpt_4056, _cvpt_4057, _cvpt_4058, _cvpt_4059, 
            _cvpt_4060, _cvpt_4061, _cvpt_4062, _cvpt_4063, _cvpt_4064, 
            _cvpt_4065, _cvpt_4066, _cvpt_4067, _cvpt_4068, _cvpt_4069, 
            _cvpt_4070, _cvpt_4071, _cvpt_4072, _cvpt_4073, _cvpt_4074, 
            _cvpt_4075, _cvpt_4076, _cvpt_4077, _cvpt_4078, _cvpt_4079, 
            _cvpt_4080, _cvpt_4081, _cvpt_4082, _cvpt_4083, _cvpt_4084, 
            _cvpt_4085, _cvpt_4086, _cvpt_4087, _cvpt_4088, _cvpt_4089, 
            _cvpt_4090, _cvpt_4091, _cvpt_4092, _cvpt_4093, _cvpt_4094, 
            _cvpt_4095, _cvpt_4096, _cvpt_4097, _cvpt_4098, _cvpt_4099, 
            _cvpt_4100, _cvpt_4101, _cvpt_4102, _cvpt_4103, _cvpt_4104, 
            _cvpt_4105, _cvpt_4106, _cvpt_4107, _cvpt_4108, _cvpt_4109, 
            _cvpt_4110, _cvpt_4111, _cvpt_4112, _cvpt_4113, _cvpt_4114, 
            _cvpt_4115, _cvpt_4116, _cvpt_4117, _cvpt_4118, _cvpt_4119, 
            _cvpt_4120, _cvpt_4121, _cvpt_4122, _cvpt_4123, _cvpt_4124, 
            _cvpt_4125, _cvpt_4126, _cvpt_4127, _cvpt_4128, _cvpt_4129, 
            _cvpt_4130, _cvpt_4131, _cvpt_4132, _cvpt_4133, _cvpt_4134, 
            _cvpt_4135, _cvpt_4136, _cvpt_4137, _cvpt_4138, _cvpt_4139, 
            _cvpt_4140, _cvpt_4141, _cvpt_4142, _cvpt_4143, _cvpt_4144, 
            _cvpt_4145, _cvpt_4146, _cvpt_4147, _cvpt_4148, _cvpt_4149, 
            _cvpt_4150, _cvpt_4151, _cvpt_4152, _cvpt_4153, _cvpt_4154, 
            _cvpt_4155, _cvpt_4156, _cvpt_4157, _cvpt_4158, _cvpt_4159, 
            _cvpt_4160, _cvpt_4161, _cvpt_4162, _cvpt_4163, _cvpt_4164, 
            _cvpt_4165, _cvpt_4166, _cvpt_4167, _cvpt_4168, _cvpt_4169, 
            _cvpt_4170, _cvpt_4171, _cvpt_4172, _cvpt_4173, _cvpt_4174, 
            _cvpt_4175, _cvpt_4176, _cvpt_4177, _cvpt_4178, _cvpt_4179, 
            _cvpt_4180, _cvpt_4181, _cvpt_4182, _cvpt_4183, _cvpt_4184, 
            _cvpt_4185, _cvpt_4186, _cvpt_4187, _cvpt_4188, _cvpt_4189, 
            _cvpt_4190, _cvpt_4191, _cvpt_4192, _cvpt_4193, _cvpt_4194, 
            _cvpt_4195, _cvpt_4196, _cvpt_4197, _cvpt_4198, _cvpt_4199, 
            _cvpt_4200, _cvpt_4201, _cvpt_4202, _cvpt_4203, _cvpt_4204, 
            _cvpt_4205, _cvpt_4206, _cvpt_4207, _cvpt_4208, _cvpt_4209, 
            _cvpt_4210, _cvpt_4211, _cvpt_4212, _cvpt_4213, _cvpt_4214, 
            _cvpt_4215, _cvpt_4216, _cvpt_4217, _cvpt_4218, _cvpt_4219, 
            _cvpt_4220, _cvpt_4221, _cvpt_4222, _cvpt_4223, _cvpt_4224, 
            _cvpt_4225, _cvpt_4226, _cvpt_4227, _cvpt_4228, _cvpt_4229, 
            _cvpt_4230, _cvpt_4231, _cvpt_4232, _cvpt_4233, _cvpt_4234, 
            _cvpt_4235, _cvpt_4236, _cvpt_4237, _cvpt_4238, _cvpt_4239, 
            _cvpt_4240, _cvpt_4241, _cvpt_4242, _cvpt_4243, _cvpt_4244, 
            _cvpt_4245, _cvpt_4246, _cvpt_4247, _cvpt_4248, _cvpt_4249, 
            _cvpt_4250, _cvpt_4251, _cvpt_4252, _cvpt_4253, _cvpt_4254, 
            _cvpt_4255, _cvpt_4256, _cvpt_4257, _cvpt_4258, _cvpt_4259, 
            _cvpt_4260, _cvpt_4261, _cvpt_4262, _cvpt_4263, _cvpt_4264, 
            _cvpt_4265, _cvpt_4266, _cvpt_4267, _cvpt_4268, _cvpt_4269, 
            _cvpt_4270, _cvpt_4271, _cvpt_4272, _cvpt_4273, _cvpt_4274, 
            _cvpt_4275, _cvpt_4276, _cvpt_4277, _cvpt_4278, _cvpt_4279, 
            _cvpt_4280, _cvpt_4281, _cvpt_4282, _cvpt_4283, _cvpt_4284, 
            _cvpt_4285, _cvpt_4286, _cvpt_4287, _cvpt_4288, _cvpt_4289, 
            _cvpt_4290, _cvpt_4291, _cvpt_4292, _cvpt_4293, _cvpt_4294, 
            _cvpt_4295, _cvpt_4296, _cvpt_4297, _cvpt_4298, _cvpt_4299, 
            _cvpt_4300, _cvpt_4301, _cvpt_4302, _cvpt_4303, _cvpt_4304, 
            _cvpt_4305, _cvpt_4306, _cvpt_4307, _cvpt_4308, _cvpt_4309, 
            _cvpt_4310, _cvpt_4311, _cvpt_4312, _cvpt_4313, _cvpt_4314, 
            _cvpt_4315, _cvpt_4316, _cvpt_4317, _cvpt_4318, _cvpt_4319, 
            _cvpt_4320, _cvpt_4321, _cvpt_4322, _cvpt_4323, _cvpt_4324, 
            _cvpt_4325, _cvpt_4326, _cvpt_4327, _cvpt_4328, _cvpt_4329, 
            _cvpt_4330, _cvpt_4331, _cvpt_4332, _cvpt_4333, _cvpt_4334, 
            _cvpt_4335, _cvpt_4336, _cvpt_4337, _cvpt_4338, _cvpt_4339, 
            _cvpt_4340, _cvpt_4341, _cvpt_4342, _cvpt_4343, _cvpt_4344, 
            _cvpt_4345, _cvpt_4346, _cvpt_4347, _cvpt_4348, _cvpt_4349, 
            _cvpt_4350, _cvpt_4351, _cvpt_4352, _cvpt_4353, _cvpt_4354, 
            _cvpt_4355, _cvpt_4356, _cvpt_4357, _cvpt_4358, _cvpt_4359, 
            _cvpt_4360, _cvpt_4361, _cvpt_4362, _cvpt_4363, _cvpt_4364, 
            _cvpt_4365, _cvpt_4366, _cvpt_4367, _cvpt_4368, _cvpt_4369, 
            _cvpt_4370, _cvpt_4371, _cvpt_4372, _cvpt_4373, _cvpt_4374, 
            _cvpt_4375, _cvpt_4376, _cvpt_4377, _cvpt_4378, _cvpt_4379, 
            _cvpt_4380, _cvpt_4381, _cvpt_4382, _cvpt_4383, _cvpt_4384, 
            _cvpt_4385, _cvpt_4386, _cvpt_4387, _cvpt_4388, _cvpt_4389, 
            _cvpt_4390, _cvpt_4391, _cvpt_4392, _cvpt_4393, _cvpt_4394, 
            _cvpt_4395, _cvpt_4396, _cvpt_4397, _cvpt_4398, _cvpt_4399, 
            _cvpt_4400, _cvpt_4401, _cvpt_4402, _cvpt_4403, _cvpt_4404, 
            _cvpt_4405, _cvpt_4406, _cvpt_4407, _cvpt_4408, _cvpt_4409, 
            _cvpt_4410, _cvpt_4411, _cvpt_4412, _cvpt_4413, _cvpt_4414, 
            _cvpt_4415, _cvpt_4416, _cvpt_4417, _cvpt_4418, _cvpt_4419, 
            _cvpt_4420, _cvpt_4421, _cvpt_4422, _cvpt_4423, _cvpt_4424, 
            _cvpt_4425, _cvpt_4426, _cvpt_4427, _cvpt_4428, _cvpt_4429, 
            _cvpt_4430, _cvpt_4431, _cvpt_4432, _cvpt_4433, _cvpt_4434, 
            _cvpt_4435, _cvpt_4436);   // oc8051_tb.v(104)
    input rst;   // oc8051_tb.v(112)
    input clk;   // oc8051_tb.v(112)
    output _cvpt_0;   // oc8051_tb.v(104)
    output _cvpt_1;   // oc8051_tb.v(104)
    output _cvpt_2;   // oc8051_tb.v(104)
    output _cvpt_3;   // oc8051_tb.v(104)
    output _cvpt_4;   // oc8051_tb.v(104)
    output _cvpt_5;   // oc8051_tb.v(104)
    output _cvpt_6;   // oc8051_tb.v(104)
    output _cvpt_7;   // oc8051_tb.v(104)
    output _cvpt_8;   // oc8051_tb.v(104)
    output _cvpt_9;   // oc8051_tb.v(104)
    output _cvpt_10;   // oc8051_tb.v(104)
    output _cvpt_11;   // oc8051_tb.v(104)
    output _cvpt_12;   // oc8051_tb.v(104)
    output _cvpt_13;   // oc8051_tb.v(104)
    output _cvpt_14;   // oc8051_tb.v(104)
    output _cvpt_15;   // oc8051_tb.v(104)
    output _cvpt_16;   // oc8051_tb.v(104)
    output _cvpt_17;   // oc8051_tb.v(104)
    output _cvpt_18;   // oc8051_tb.v(104)
    output _cvpt_19;   // oc8051_tb.v(104)
    output _cvpt_20;   // oc8051_tb.v(104)
    output _cvpt_21;   // oc8051_tb.v(104)
    output _cvpt_22;   // oc8051_tb.v(104)
    output _cvpt_23;   // oc8051_tb.v(104)
    output _cvpt_24;   // oc8051_tb.v(104)
    output _cvpt_25;   // oc8051_tb.v(104)
    output _cvpt_26;   // oc8051_tb.v(104)
    output _cvpt_27;   // oc8051_tb.v(104)
    output _cvpt_28;   // oc8051_tb.v(104)
    output _cvpt_29;   // oc8051_tb.v(104)
    output _cvpt_30;   // oc8051_tb.v(104)
    output _cvpt_31;   // oc8051_tb.v(104)
    output _cvpt_32;   // oc8051_tb.v(104)
    output _cvpt_33;   // oc8051_tb.v(104)
    output _cvpt_34;   // oc8051_tb.v(104)
    output _cvpt_35;   // oc8051_tb.v(104)
    output _cvpt_36;   // oc8051_tb.v(104)
    output _cvpt_37;   // oc8051_tb.v(104)
    output _cvpt_38;   // oc8051_tb.v(104)
    output _cvpt_39;   // oc8051_tb.v(104)
    output _cvpt_40;   // oc8051_tb.v(104)
    output _cvpt_41;   // oc8051_tb.v(104)
    output _cvpt_42;   // oc8051_tb.v(104)
    output _cvpt_43;   // oc8051_tb.v(104)
    output _cvpt_44;   // oc8051_tb.v(104)
    output _cvpt_45;   // oc8051_tb.v(104)
    output _cvpt_46;   // oc8051_tb.v(104)
    output _cvpt_47;   // oc8051_tb.v(104)
    output _cvpt_48;   // oc8051_tb.v(104)
    output _cvpt_49;   // oc8051_tb.v(104)
    output _cvpt_50;   // oc8051_tb.v(104)
    output _cvpt_51;   // oc8051_tb.v(104)
    output _cvpt_52;   // oc8051_tb.v(104)
    output _cvpt_53;   // oc8051_tb.v(104)
    output _cvpt_54;   // oc8051_tb.v(104)
    output _cvpt_55;   // oc8051_tb.v(104)
    output _cvpt_56;   // oc8051_tb.v(104)
    output _cvpt_57;   // oc8051_tb.v(104)
    output _cvpt_58;   // oc8051_tb.v(104)
    output _cvpt_59;   // oc8051_tb.v(104)
    output _cvpt_60;   // oc8051_tb.v(104)
    output _cvpt_61;   // oc8051_tb.v(104)
    output _cvpt_62;   // oc8051_tb.v(104)
    output _cvpt_63;   // oc8051_tb.v(104)
    output _cvpt_64;   // oc8051_tb.v(104)
    output _cvpt_65;   // oc8051_tb.v(104)
    output _cvpt_66;   // oc8051_tb.v(104)
    output _cvpt_67;   // oc8051_tb.v(104)
    output _cvpt_68;   // oc8051_tb.v(104)
    output _cvpt_69;   // oc8051_tb.v(104)
    output _cvpt_70;   // oc8051_tb.v(104)
    output _cvpt_71;   // oc8051_tb.v(104)
    output _cvpt_72;   // oc8051_tb.v(104)
    output _cvpt_73;   // oc8051_tb.v(104)
    output _cvpt_74;   // oc8051_tb.v(104)
    output _cvpt_75;   // oc8051_tb.v(104)
    output _cvpt_76;   // oc8051_tb.v(104)
    output _cvpt_77;   // oc8051_tb.v(104)
    output _cvpt_78;   // oc8051_tb.v(104)
    output _cvpt_79;   // oc8051_tb.v(104)
    output _cvpt_80;   // oc8051_tb.v(104)
    output _cvpt_81;   // oc8051_tb.v(104)
    output _cvpt_82;   // oc8051_tb.v(104)
    output _cvpt_83;   // oc8051_tb.v(104)
    output _cvpt_84;   // oc8051_tb.v(104)
    output _cvpt_85;   // oc8051_tb.v(104)
    output _cvpt_86;   // oc8051_tb.v(104)
    output _cvpt_87;   // oc8051_tb.v(104)
    output _cvpt_88;   // oc8051_tb.v(104)
    output _cvpt_89;   // oc8051_tb.v(104)
    output _cvpt_90;   // oc8051_tb.v(104)
    output _cvpt_91;   // oc8051_tb.v(104)
    output _cvpt_92;   // oc8051_tb.v(104)
    output _cvpt_93;   // oc8051_tb.v(104)
    output _cvpt_94;   // oc8051_tb.v(104)
    output _cvpt_95;   // oc8051_tb.v(104)
    output _cvpt_96;   // oc8051_tb.v(104)
    output _cvpt_97;   // oc8051_tb.v(104)
    output _cvpt_98;   // oc8051_tb.v(104)
    output _cvpt_99;   // oc8051_tb.v(104)
    output _cvpt_100;   // oc8051_tb.v(104)
    output _cvpt_101;   // oc8051_tb.v(104)
    output _cvpt_102;   // oc8051_tb.v(104)
    output _cvpt_103;   // oc8051_tb.v(104)
    output _cvpt_104;   // oc8051_tb.v(104)
    output _cvpt_105;   // oc8051_tb.v(104)
    output _cvpt_106;   // oc8051_tb.v(104)
    output _cvpt_107;   // oc8051_tb.v(104)
    output _cvpt_108;   // oc8051_tb.v(104)
    output _cvpt_109;   // oc8051_tb.v(104)
    output _cvpt_110;   // oc8051_tb.v(104)
    output _cvpt_111;   // oc8051_tb.v(104)
    output _cvpt_112;   // oc8051_tb.v(104)
    output _cvpt_113;   // oc8051_tb.v(104)
    output _cvpt_114;   // oc8051_tb.v(104)
    output _cvpt_115;   // oc8051_tb.v(104)
    output _cvpt_116;   // oc8051_tb.v(104)
    output _cvpt_117;   // oc8051_tb.v(104)
    output _cvpt_118;   // oc8051_tb.v(104)
    output _cvpt_119;   // oc8051_tb.v(104)
    output _cvpt_120;   // oc8051_tb.v(104)
    output _cvpt_121;   // oc8051_tb.v(104)
    output _cvpt_122;   // oc8051_tb.v(104)
    output _cvpt_123;   // oc8051_tb.v(104)
    output _cvpt_124;   // oc8051_tb.v(104)
    output _cvpt_125;   // oc8051_tb.v(104)
    output _cvpt_126;   // oc8051_tb.v(104)
    output _cvpt_127;   // oc8051_tb.v(104)
    output _cvpt_128;   // oc8051_tb.v(104)
    output _cvpt_129;   // oc8051_tb.v(104)
    output _cvpt_130;   // oc8051_tb.v(104)
    output _cvpt_131;   // oc8051_tb.v(104)
    output _cvpt_132;   // oc8051_tb.v(104)
    output _cvpt_133;   // oc8051_tb.v(104)
    output _cvpt_134;   // oc8051_tb.v(104)
    output _cvpt_135;   // oc8051_tb.v(104)
    output _cvpt_136;   // oc8051_tb.v(104)
    output _cvpt_137;   // oc8051_tb.v(104)
    output _cvpt_138;   // oc8051_tb.v(104)
    output _cvpt_139;   // oc8051_tb.v(104)
    output _cvpt_140;   // oc8051_tb.v(104)
    output _cvpt_141;   // oc8051_tb.v(104)
    output _cvpt_142;   // oc8051_tb.v(104)
    output _cvpt_143;   // oc8051_tb.v(104)
    output _cvpt_144;   // oc8051_tb.v(104)
    output _cvpt_145;   // oc8051_tb.v(104)
    output _cvpt_146;   // oc8051_tb.v(104)
    output _cvpt_147;   // oc8051_tb.v(104)
    output _cvpt_148;   // oc8051_tb.v(104)
    output _cvpt_149;   // oc8051_tb.v(104)
    output _cvpt_150;   // oc8051_tb.v(104)
    output _cvpt_151;   // oc8051_tb.v(104)
    output _cvpt_152;   // oc8051_tb.v(104)
    output _cvpt_153;   // oc8051_tb.v(104)
    output _cvpt_154;   // oc8051_tb.v(104)
    output _cvpt_155;   // oc8051_tb.v(104)
    output _cvpt_156;   // oc8051_tb.v(104)
    output _cvpt_157;   // oc8051_tb.v(104)
    output _cvpt_158;   // oc8051_tb.v(104)
    output _cvpt_159;   // oc8051_tb.v(104)
    output _cvpt_160;   // oc8051_tb.v(104)
    output _cvpt_161;   // oc8051_tb.v(104)
    output _cvpt_162;   // oc8051_tb.v(104)
    output _cvpt_163;   // oc8051_tb.v(104)
    output _cvpt_164;   // oc8051_tb.v(104)
    output _cvpt_165;   // oc8051_tb.v(104)
    output _cvpt_166;   // oc8051_tb.v(104)
    output _cvpt_167;   // oc8051_tb.v(104)
    output _cvpt_168;   // oc8051_tb.v(104)
    output _cvpt_169;   // oc8051_tb.v(104)
    output _cvpt_170;   // oc8051_tb.v(104)
    output _cvpt_171;   // oc8051_tb.v(104)
    output _cvpt_172;   // oc8051_tb.v(104)
    output _cvpt_173;   // oc8051_tb.v(104)
    output _cvpt_174;   // oc8051_tb.v(104)
    output _cvpt_175;   // oc8051_tb.v(104)
    output _cvpt_176;   // oc8051_tb.v(104)
    output _cvpt_177;   // oc8051_tb.v(104)
    output _cvpt_178;   // oc8051_tb.v(104)
    output _cvpt_179;   // oc8051_tb.v(104)
    output _cvpt_180;   // oc8051_tb.v(104)
    output _cvpt_181;   // oc8051_tb.v(104)
    output _cvpt_182;   // oc8051_tb.v(104)
    output _cvpt_183;   // oc8051_tb.v(104)
    output _cvpt_184;   // oc8051_tb.v(104)
    output _cvpt_185;   // oc8051_tb.v(104)
    output _cvpt_186;   // oc8051_tb.v(104)
    output _cvpt_187;   // oc8051_tb.v(104)
    output _cvpt_188;   // oc8051_tb.v(104)
    output _cvpt_189;   // oc8051_tb.v(104)
    output _cvpt_190;   // oc8051_tb.v(104)
    output _cvpt_191;   // oc8051_tb.v(104)
    output _cvpt_192;   // oc8051_tb.v(104)
    output _cvpt_193;   // oc8051_tb.v(104)
    output _cvpt_194;   // oc8051_tb.v(104)
    output _cvpt_195;   // oc8051_tb.v(104)
    output _cvpt_196;   // oc8051_tb.v(104)
    output _cvpt_197;   // oc8051_tb.v(104)
    output _cvpt_198;   // oc8051_tb.v(104)
    output _cvpt_199;   // oc8051_tb.v(104)
    output _cvpt_200;   // oc8051_tb.v(104)
    output _cvpt_201;   // oc8051_tb.v(104)
    output _cvpt_202;   // oc8051_tb.v(104)
    output _cvpt_203;   // oc8051_tb.v(104)
    output _cvpt_204;   // oc8051_tb.v(104)
    output _cvpt_205;   // oc8051_tb.v(104)
    output _cvpt_206;   // oc8051_tb.v(104)
    output _cvpt_207;   // oc8051_tb.v(104)
    output _cvpt_208;   // oc8051_tb.v(104)
    output _cvpt_209;   // oc8051_tb.v(104)
    output _cvpt_210;   // oc8051_tb.v(104)
    output _cvpt_211;   // oc8051_tb.v(104)
    output _cvpt_212;   // oc8051_tb.v(104)
    output _cvpt_213;   // oc8051_tb.v(104)
    output _cvpt_214;   // oc8051_tb.v(104)
    output _cvpt_215;   // oc8051_tb.v(104)
    output _cvpt_216;   // oc8051_tb.v(104)
    output _cvpt_217;   // oc8051_tb.v(104)
    output _cvpt_218;   // oc8051_tb.v(104)
    output _cvpt_219;   // oc8051_tb.v(104)
    output _cvpt_220;   // oc8051_tb.v(104)
    output _cvpt_221;   // oc8051_tb.v(104)
    output _cvpt_222;   // oc8051_tb.v(104)
    output _cvpt_223;   // oc8051_tb.v(104)
    output _cvpt_224;   // oc8051_tb.v(104)
    output _cvpt_225;   // oc8051_tb.v(104)
    output _cvpt_226;   // oc8051_tb.v(104)
    output _cvpt_227;   // oc8051_tb.v(104)
    output _cvpt_228;   // oc8051_tb.v(104)
    output _cvpt_229;   // oc8051_tb.v(104)
    output _cvpt_230;   // oc8051_tb.v(104)
    output _cvpt_231;   // oc8051_tb.v(104)
    output _cvpt_232;   // oc8051_tb.v(104)
    output _cvpt_233;   // oc8051_tb.v(104)
    output _cvpt_234;   // oc8051_tb.v(104)
    output _cvpt_235;   // oc8051_tb.v(104)
    output _cvpt_236;   // oc8051_tb.v(104)
    output _cvpt_237;   // oc8051_tb.v(104)
    output _cvpt_238;   // oc8051_tb.v(104)
    output _cvpt_239;   // oc8051_tb.v(104)
    output _cvpt_240;   // oc8051_tb.v(104)
    output _cvpt_241;   // oc8051_tb.v(104)
    output _cvpt_242;   // oc8051_tb.v(104)
    output _cvpt_243;   // oc8051_tb.v(104)
    output _cvpt_244;   // oc8051_tb.v(104)
    output _cvpt_245;   // oc8051_tb.v(104)
    output _cvpt_246;   // oc8051_tb.v(104)
    output _cvpt_247;   // oc8051_tb.v(104)
    output _cvpt_248;   // oc8051_tb.v(104)
    output _cvpt_249;   // oc8051_tb.v(104)
    output _cvpt_250;   // oc8051_tb.v(104)
    output _cvpt_251;   // oc8051_tb.v(104)
    output _cvpt_252;   // oc8051_tb.v(104)
    output _cvpt_253;   // oc8051_tb.v(104)
    output _cvpt_254;   // oc8051_tb.v(104)
    output _cvpt_255;   // oc8051_tb.v(104)
    output _cvpt_256;   // oc8051_tb.v(104)
    output _cvpt_257;   // oc8051_tb.v(104)
    output _cvpt_258;   // oc8051_tb.v(104)
    output _cvpt_259;   // oc8051_tb.v(104)
    output _cvpt_260;   // oc8051_tb.v(104)
    output _cvpt_261;   // oc8051_tb.v(104)
    output _cvpt_262;   // oc8051_tb.v(104)
    output _cvpt_263;   // oc8051_tb.v(104)
    output _cvpt_264;   // oc8051_tb.v(104)
    output _cvpt_265;   // oc8051_tb.v(104)
    output _cvpt_266;   // oc8051_tb.v(104)
    output _cvpt_267;   // oc8051_tb.v(104)
    output _cvpt_268;   // oc8051_tb.v(104)
    output _cvpt_269;   // oc8051_tb.v(104)
    output _cvpt_270;   // oc8051_tb.v(104)
    output _cvpt_271;   // oc8051_tb.v(104)
    output _cvpt_272;   // oc8051_tb.v(104)
    output _cvpt_273;   // oc8051_tb.v(104)
    output _cvpt_274;   // oc8051_tb.v(104)
    output _cvpt_275;   // oc8051_tb.v(104)
    output _cvpt_276;   // oc8051_tb.v(104)
    output _cvpt_277;   // oc8051_tb.v(104)
    output _cvpt_278;   // oc8051_tb.v(104)
    output _cvpt_279;   // oc8051_tb.v(104)
    output _cvpt_280;   // oc8051_tb.v(104)
    output _cvpt_281;   // oc8051_tb.v(104)
    output _cvpt_282;   // oc8051_tb.v(104)
    output _cvpt_283;   // oc8051_tb.v(104)
    output _cvpt_284;   // oc8051_tb.v(104)
    output _cvpt_285;   // oc8051_tb.v(104)
    output _cvpt_286;   // oc8051_tb.v(104)
    output _cvpt_287;   // oc8051_tb.v(104)
    output _cvpt_288;   // oc8051_tb.v(104)
    output _cvpt_289;   // oc8051_tb.v(104)
    output _cvpt_290;   // oc8051_tb.v(104)
    output _cvpt_291;   // oc8051_tb.v(104)
    output _cvpt_292;   // oc8051_tb.v(104)
    output _cvpt_293;   // oc8051_tb.v(104)
    output _cvpt_294;   // oc8051_tb.v(104)
    output _cvpt_295;   // oc8051_tb.v(104)
    output _cvpt_296;   // oc8051_tb.v(104)
    output _cvpt_297;   // oc8051_tb.v(104)
    output _cvpt_298;   // oc8051_tb.v(104)
    output _cvpt_299;   // oc8051_tb.v(104)
    output _cvpt_300;   // oc8051_tb.v(104)
    output _cvpt_301;   // oc8051_tb.v(104)
    output _cvpt_302;   // oc8051_tb.v(104)
    output _cvpt_303;   // oc8051_tb.v(104)
    output _cvpt_304;   // oc8051_tb.v(104)
    output _cvpt_305;   // oc8051_tb.v(104)
    output _cvpt_306;   // oc8051_tb.v(104)
    output _cvpt_307;   // oc8051_tb.v(104)
    output _cvpt_308;   // oc8051_tb.v(104)
    output _cvpt_309;   // oc8051_tb.v(104)
    output _cvpt_310;   // oc8051_tb.v(104)
    output _cvpt_311;   // oc8051_tb.v(104)
    output _cvpt_312;   // oc8051_tb.v(104)
    output _cvpt_313;   // oc8051_tb.v(104)
    output _cvpt_314;   // oc8051_tb.v(104)
    output _cvpt_315;   // oc8051_tb.v(104)
    output _cvpt_316;   // oc8051_tb.v(104)
    output _cvpt_317;   // oc8051_tb.v(104)
    output _cvpt_318;   // oc8051_tb.v(104)
    output _cvpt_319;   // oc8051_tb.v(104)
    output _cvpt_320;   // oc8051_tb.v(104)
    output _cvpt_321;   // oc8051_tb.v(104)
    output _cvpt_322;   // oc8051_tb.v(104)
    output _cvpt_323;   // oc8051_tb.v(104)
    output _cvpt_324;   // oc8051_tb.v(104)
    output _cvpt_325;   // oc8051_tb.v(104)
    output _cvpt_326;   // oc8051_tb.v(104)
    output _cvpt_327;   // oc8051_tb.v(104)
    output _cvpt_328;   // oc8051_tb.v(104)
    output _cvpt_329;   // oc8051_tb.v(104)
    output _cvpt_330;   // oc8051_tb.v(104)
    output _cvpt_331;   // oc8051_tb.v(104)
    output _cvpt_332;   // oc8051_tb.v(104)
    output _cvpt_333;   // oc8051_tb.v(104)
    output _cvpt_334;   // oc8051_tb.v(104)
    output _cvpt_335;   // oc8051_tb.v(104)
    output _cvpt_336;   // oc8051_tb.v(104)
    output _cvpt_337;   // oc8051_tb.v(104)
    output _cvpt_338;   // oc8051_tb.v(104)
    output _cvpt_339;   // oc8051_tb.v(104)
    output _cvpt_340;   // oc8051_tb.v(104)
    output _cvpt_341;   // oc8051_tb.v(104)
    output _cvpt_342;   // oc8051_tb.v(104)
    output _cvpt_343;   // oc8051_tb.v(104)
    output _cvpt_344;   // oc8051_tb.v(104)
    output _cvpt_345;   // oc8051_tb.v(104)
    output _cvpt_346;   // oc8051_tb.v(104)
    output _cvpt_347;   // oc8051_tb.v(104)
    output _cvpt_348;   // oc8051_tb.v(104)
    output _cvpt_349;   // oc8051_tb.v(104)
    output _cvpt_350;   // oc8051_tb.v(104)
    output _cvpt_351;   // oc8051_tb.v(104)
    output _cvpt_352;   // oc8051_tb.v(104)
    output _cvpt_353;   // oc8051_tb.v(104)
    output _cvpt_354;   // oc8051_tb.v(104)
    output _cvpt_355;   // oc8051_tb.v(104)
    output _cvpt_356;   // oc8051_tb.v(104)
    output _cvpt_357;   // oc8051_tb.v(104)
    output _cvpt_358;   // oc8051_tb.v(104)
    output _cvpt_359;   // oc8051_tb.v(104)
    output _cvpt_360;   // oc8051_tb.v(104)
    output _cvpt_361;   // oc8051_tb.v(104)
    output _cvpt_362;   // oc8051_tb.v(104)
    output _cvpt_363;   // oc8051_tb.v(104)
    output _cvpt_364;   // oc8051_tb.v(104)
    output _cvpt_365;   // oc8051_tb.v(104)
    output _cvpt_366;   // oc8051_tb.v(104)
    output _cvpt_367;   // oc8051_tb.v(104)
    output _cvpt_368;   // oc8051_tb.v(104)
    output _cvpt_369;   // oc8051_tb.v(104)
    output _cvpt_370;   // oc8051_tb.v(104)
    output _cvpt_371;   // oc8051_tb.v(104)
    output _cvpt_372;   // oc8051_tb.v(104)
    output _cvpt_373;   // oc8051_tb.v(104)
    output _cvpt_374;   // oc8051_tb.v(104)
    output _cvpt_375;   // oc8051_tb.v(104)
    output _cvpt_376;   // oc8051_tb.v(104)
    output _cvpt_377;   // oc8051_tb.v(104)
    output _cvpt_378;   // oc8051_tb.v(104)
    output _cvpt_379;   // oc8051_tb.v(104)
    output _cvpt_380;   // oc8051_tb.v(104)
    output _cvpt_381;   // oc8051_tb.v(104)
    output _cvpt_382;   // oc8051_tb.v(104)
    output _cvpt_383;   // oc8051_tb.v(104)
    output _cvpt_384;   // oc8051_tb.v(104)
    output _cvpt_385;   // oc8051_tb.v(104)
    output _cvpt_386;   // oc8051_tb.v(104)
    output _cvpt_387;   // oc8051_tb.v(104)
    output _cvpt_388;   // oc8051_tb.v(104)
    output _cvpt_389;   // oc8051_tb.v(104)
    output _cvpt_390;   // oc8051_tb.v(104)
    output _cvpt_391;   // oc8051_tb.v(104)
    output _cvpt_392;   // oc8051_tb.v(104)
    output _cvpt_393;   // oc8051_tb.v(104)
    output _cvpt_394;   // oc8051_tb.v(104)
    output _cvpt_395;   // oc8051_tb.v(104)
    output _cvpt_396;   // oc8051_tb.v(104)
    output _cvpt_397;   // oc8051_tb.v(104)
    output _cvpt_398;   // oc8051_tb.v(104)
    output _cvpt_399;   // oc8051_tb.v(104)
    output _cvpt_400;   // oc8051_tb.v(104)
    output _cvpt_401;   // oc8051_tb.v(104)
    output _cvpt_402;   // oc8051_tb.v(104)
    output _cvpt_403;   // oc8051_tb.v(104)
    output _cvpt_404;   // oc8051_tb.v(104)
    output _cvpt_405;   // oc8051_tb.v(104)
    output _cvpt_406;   // oc8051_tb.v(104)
    output _cvpt_407;   // oc8051_tb.v(104)
    output _cvpt_408;   // oc8051_tb.v(104)
    output _cvpt_409;   // oc8051_tb.v(104)
    output _cvpt_410;   // oc8051_tb.v(104)
    output _cvpt_411;   // oc8051_tb.v(104)
    output _cvpt_412;   // oc8051_tb.v(104)
    output _cvpt_413;   // oc8051_tb.v(104)
    output _cvpt_414;   // oc8051_tb.v(104)
    output _cvpt_415;   // oc8051_tb.v(104)
    output _cvpt_416;   // oc8051_tb.v(104)
    output _cvpt_417;   // oc8051_tb.v(104)
    output _cvpt_418;   // oc8051_tb.v(104)
    output _cvpt_419;   // oc8051_tb.v(104)
    output _cvpt_420;   // oc8051_tb.v(104)
    output _cvpt_421;   // oc8051_tb.v(104)
    output _cvpt_422;   // oc8051_tb.v(104)
    output _cvpt_423;   // oc8051_tb.v(104)
    output _cvpt_424;   // oc8051_tb.v(104)
    output _cvpt_425;   // oc8051_tb.v(104)
    output _cvpt_426;   // oc8051_tb.v(104)
    output _cvpt_427;   // oc8051_tb.v(104)
    output _cvpt_428;   // oc8051_tb.v(104)
    output _cvpt_429;   // oc8051_tb.v(104)
    output _cvpt_430;   // oc8051_tb.v(104)
    output _cvpt_431;   // oc8051_tb.v(104)
    output _cvpt_432;   // oc8051_tb.v(104)
    output _cvpt_433;   // oc8051_tb.v(104)
    output _cvpt_434;   // oc8051_tb.v(104)
    output _cvpt_435;   // oc8051_tb.v(104)
    output _cvpt_436;   // oc8051_tb.v(104)
    output _cvpt_437;   // oc8051_tb.v(104)
    output _cvpt_438;   // oc8051_tb.v(104)
    output _cvpt_439;   // oc8051_tb.v(104)
    output _cvpt_440;   // oc8051_tb.v(104)
    output _cvpt_441;   // oc8051_tb.v(104)
    output _cvpt_442;   // oc8051_tb.v(104)
    output _cvpt_443;   // oc8051_tb.v(104)
    output _cvpt_444;   // oc8051_tb.v(104)
    output _cvpt_445;   // oc8051_tb.v(104)
    output _cvpt_446;   // oc8051_tb.v(104)
    output _cvpt_447;   // oc8051_tb.v(104)
    output _cvpt_448;   // oc8051_tb.v(104)
    output _cvpt_449;   // oc8051_tb.v(104)
    output _cvpt_450;   // oc8051_tb.v(104)
    output _cvpt_451;   // oc8051_tb.v(104)
    output _cvpt_452;   // oc8051_tb.v(104)
    output _cvpt_453;   // oc8051_tb.v(104)
    output _cvpt_454;   // oc8051_tb.v(104)
    output _cvpt_455;   // oc8051_tb.v(104)
    output _cvpt_456;   // oc8051_tb.v(104)
    output _cvpt_457;   // oc8051_tb.v(104)
    output _cvpt_458;   // oc8051_tb.v(104)
    output _cvpt_459;   // oc8051_tb.v(104)
    output _cvpt_460;   // oc8051_tb.v(104)
    output _cvpt_461;   // oc8051_tb.v(104)
    output _cvpt_462;   // oc8051_tb.v(104)
    output _cvpt_463;   // oc8051_tb.v(104)
    output _cvpt_464;   // oc8051_tb.v(104)
    output _cvpt_465;   // oc8051_tb.v(104)
    output _cvpt_466;   // oc8051_tb.v(104)
    output _cvpt_467;   // oc8051_tb.v(104)
    output _cvpt_468;   // oc8051_tb.v(104)
    output _cvpt_469;   // oc8051_tb.v(104)
    output _cvpt_470;   // oc8051_tb.v(104)
    output _cvpt_471;   // oc8051_tb.v(104)
    output _cvpt_472;   // oc8051_tb.v(104)
    output _cvpt_473;   // oc8051_tb.v(104)
    output _cvpt_474;   // oc8051_tb.v(104)
    output _cvpt_475;   // oc8051_tb.v(104)
    output _cvpt_476;   // oc8051_tb.v(104)
    output _cvpt_477;   // oc8051_tb.v(104)
    output _cvpt_478;   // oc8051_tb.v(104)
    output _cvpt_479;   // oc8051_tb.v(104)
    output _cvpt_480;   // oc8051_tb.v(104)
    output _cvpt_481;   // oc8051_tb.v(104)
    output _cvpt_482;   // oc8051_tb.v(104)
    output _cvpt_483;   // oc8051_tb.v(104)
    output _cvpt_484;   // oc8051_tb.v(104)
    output _cvpt_485;   // oc8051_tb.v(104)
    output _cvpt_486;   // oc8051_tb.v(104)
    output _cvpt_487;   // oc8051_tb.v(104)
    output _cvpt_488;   // oc8051_tb.v(104)
    output _cvpt_489;   // oc8051_tb.v(104)
    output _cvpt_490;   // oc8051_tb.v(104)
    output _cvpt_491;   // oc8051_tb.v(104)
    output _cvpt_492;   // oc8051_tb.v(104)
    output _cvpt_493;   // oc8051_tb.v(104)
    output _cvpt_494;   // oc8051_tb.v(104)
    output _cvpt_495;   // oc8051_tb.v(104)
    output _cvpt_496;   // oc8051_tb.v(104)
    output _cvpt_497;   // oc8051_tb.v(104)
    output _cvpt_498;   // oc8051_tb.v(104)
    output _cvpt_499;   // oc8051_tb.v(104)
    output _cvpt_500;   // oc8051_tb.v(104)
    output _cvpt_501;   // oc8051_tb.v(104)
    output _cvpt_502;   // oc8051_tb.v(104)
    output _cvpt_503;   // oc8051_tb.v(104)
    output _cvpt_504;   // oc8051_tb.v(104)
    output _cvpt_505;   // oc8051_tb.v(104)
    output _cvpt_506;   // oc8051_tb.v(104)
    output _cvpt_507;   // oc8051_tb.v(104)
    output _cvpt_508;   // oc8051_tb.v(104)
    output _cvpt_509;   // oc8051_tb.v(104)
    output _cvpt_510;   // oc8051_tb.v(104)
    output _cvpt_511;   // oc8051_tb.v(104)
    output _cvpt_512;   // oc8051_tb.v(104)
    output _cvpt_513;   // oc8051_tb.v(104)
    output _cvpt_514;   // oc8051_tb.v(104)
    output _cvpt_515;   // oc8051_tb.v(104)
    output _cvpt_516;   // oc8051_tb.v(104)
    output _cvpt_517;   // oc8051_tb.v(104)
    output _cvpt_518;   // oc8051_tb.v(104)
    output _cvpt_519;   // oc8051_tb.v(104)
    output _cvpt_520;   // oc8051_tb.v(104)
    output _cvpt_521;   // oc8051_tb.v(104)
    output _cvpt_522;   // oc8051_tb.v(104)
    output _cvpt_523;   // oc8051_tb.v(104)
    output _cvpt_524;   // oc8051_tb.v(104)
    output _cvpt_525;   // oc8051_tb.v(104)
    output _cvpt_526;   // oc8051_tb.v(104)
    output _cvpt_527;   // oc8051_tb.v(104)
    output _cvpt_528;   // oc8051_tb.v(104)
    output _cvpt_529;   // oc8051_tb.v(104)
    output _cvpt_530;   // oc8051_tb.v(104)
    output _cvpt_531;   // oc8051_tb.v(104)
    output _cvpt_532;   // oc8051_tb.v(104)
    output _cvpt_533;   // oc8051_tb.v(104)
    output _cvpt_534;   // oc8051_tb.v(104)
    output _cvpt_535;   // oc8051_tb.v(104)
    output _cvpt_536;   // oc8051_tb.v(104)
    output _cvpt_537;   // oc8051_tb.v(104)
    output _cvpt_538;   // oc8051_tb.v(104)
    output _cvpt_539;   // oc8051_tb.v(104)
    output _cvpt_540;   // oc8051_tb.v(104)
    output _cvpt_541;   // oc8051_tb.v(104)
    output _cvpt_542;   // oc8051_tb.v(104)
    output _cvpt_543;   // oc8051_tb.v(104)
    output _cvpt_544;   // oc8051_tb.v(104)
    output _cvpt_545;   // oc8051_tb.v(104)
    output _cvpt_546;   // oc8051_tb.v(104)
    output _cvpt_547;   // oc8051_tb.v(104)
    output _cvpt_548;   // oc8051_tb.v(104)
    output _cvpt_549;   // oc8051_tb.v(104)
    output _cvpt_550;   // oc8051_tb.v(104)
    output _cvpt_551;   // oc8051_tb.v(104)
    output _cvpt_552;   // oc8051_tb.v(104)
    output _cvpt_553;   // oc8051_tb.v(104)
    output _cvpt_554;   // oc8051_tb.v(104)
    output _cvpt_555;   // oc8051_tb.v(104)
    output _cvpt_556;   // oc8051_tb.v(104)
    output _cvpt_557;   // oc8051_tb.v(104)
    output _cvpt_558;   // oc8051_tb.v(104)
    output _cvpt_559;   // oc8051_tb.v(104)
    output _cvpt_560;   // oc8051_tb.v(104)
    output _cvpt_561;   // oc8051_tb.v(104)
    output _cvpt_562;   // oc8051_tb.v(104)
    output _cvpt_563;   // oc8051_tb.v(104)
    output _cvpt_564;   // oc8051_tb.v(104)
    output _cvpt_565;   // oc8051_tb.v(104)
    output _cvpt_566;   // oc8051_tb.v(104)
    output _cvpt_567;   // oc8051_tb.v(104)
    output _cvpt_568;   // oc8051_tb.v(104)
    output _cvpt_569;   // oc8051_tb.v(104)
    output _cvpt_570;   // oc8051_tb.v(104)
    output _cvpt_571;   // oc8051_tb.v(104)
    output _cvpt_572;   // oc8051_tb.v(104)
    output _cvpt_573;   // oc8051_tb.v(104)
    output _cvpt_574;   // oc8051_tb.v(104)
    output _cvpt_575;   // oc8051_tb.v(104)
    output _cvpt_576;   // oc8051_tb.v(104)
    output _cvpt_577;   // oc8051_tb.v(104)
    output _cvpt_578;   // oc8051_tb.v(104)
    output _cvpt_579;   // oc8051_tb.v(104)
    output _cvpt_580;   // oc8051_tb.v(104)
    output _cvpt_581;   // oc8051_tb.v(104)
    output _cvpt_582;   // oc8051_tb.v(104)
    output _cvpt_583;   // oc8051_tb.v(104)
    output _cvpt_584;   // oc8051_tb.v(104)
    output _cvpt_585;   // oc8051_tb.v(104)
    output _cvpt_586;   // oc8051_tb.v(104)
    output _cvpt_587;   // oc8051_tb.v(104)
    output _cvpt_588;   // oc8051_tb.v(104)
    output _cvpt_589;   // oc8051_tb.v(104)
    output _cvpt_590;   // oc8051_tb.v(104)
    output _cvpt_591;   // oc8051_tb.v(104)
    output _cvpt_592;   // oc8051_tb.v(104)
    output _cvpt_593;   // oc8051_tb.v(104)
    output _cvpt_594;   // oc8051_tb.v(104)
    output _cvpt_595;   // oc8051_tb.v(104)
    output _cvpt_596;   // oc8051_tb.v(104)
    output _cvpt_597;   // oc8051_tb.v(104)
    output _cvpt_598;   // oc8051_tb.v(104)
    output _cvpt_599;   // oc8051_tb.v(104)
    output _cvpt_600;   // oc8051_tb.v(104)
    output _cvpt_601;   // oc8051_tb.v(104)
    output _cvpt_602;   // oc8051_tb.v(104)
    output _cvpt_603;   // oc8051_tb.v(104)
    output _cvpt_604;   // oc8051_tb.v(104)
    output _cvpt_605;   // oc8051_tb.v(104)
    output _cvpt_606;   // oc8051_tb.v(104)
    output _cvpt_607;   // oc8051_tb.v(104)
    output _cvpt_608;   // oc8051_tb.v(104)
    output _cvpt_609;   // oc8051_tb.v(104)
    output _cvpt_610;   // oc8051_tb.v(104)
    output _cvpt_611;   // oc8051_tb.v(104)
    output _cvpt_612;   // oc8051_tb.v(104)
    output _cvpt_613;   // oc8051_tb.v(104)
    output _cvpt_614;   // oc8051_tb.v(104)
    output _cvpt_615;   // oc8051_tb.v(104)
    output _cvpt_616;   // oc8051_tb.v(104)
    output _cvpt_617;   // oc8051_tb.v(104)
    output _cvpt_618;   // oc8051_tb.v(104)
    output _cvpt_619;   // oc8051_tb.v(104)
    output _cvpt_620;   // oc8051_tb.v(104)
    output _cvpt_621;   // oc8051_tb.v(104)
    output _cvpt_622;   // oc8051_tb.v(104)
    output _cvpt_623;   // oc8051_tb.v(104)
    output _cvpt_624;   // oc8051_tb.v(104)
    output _cvpt_625;   // oc8051_tb.v(104)
    output _cvpt_626;   // oc8051_tb.v(104)
    output _cvpt_627;   // oc8051_tb.v(104)
    output _cvpt_628;   // oc8051_tb.v(104)
    output _cvpt_629;   // oc8051_tb.v(104)
    output _cvpt_630;   // oc8051_tb.v(104)
    output _cvpt_631;   // oc8051_tb.v(104)
    output _cvpt_632;   // oc8051_tb.v(104)
    output _cvpt_633;   // oc8051_tb.v(104)
    output _cvpt_634;   // oc8051_tb.v(104)
    output _cvpt_635;   // oc8051_tb.v(104)
    output _cvpt_636;   // oc8051_tb.v(104)
    output _cvpt_637;   // oc8051_tb.v(104)
    output _cvpt_638;   // oc8051_tb.v(104)
    output _cvpt_639;   // oc8051_tb.v(104)
    output _cvpt_640;   // oc8051_tb.v(104)
    output _cvpt_641;   // oc8051_tb.v(104)
    output _cvpt_642;   // oc8051_tb.v(104)
    output _cvpt_643;   // oc8051_tb.v(104)
    output _cvpt_644;   // oc8051_tb.v(104)
    output _cvpt_645;   // oc8051_tb.v(104)
    output _cvpt_646;   // oc8051_tb.v(104)
    output _cvpt_647;   // oc8051_tb.v(104)
    output _cvpt_648;   // oc8051_tb.v(104)
    output _cvpt_649;   // oc8051_tb.v(104)
    output _cvpt_650;   // oc8051_tb.v(104)
    output _cvpt_651;   // oc8051_tb.v(104)
    output _cvpt_652;   // oc8051_tb.v(104)
    output _cvpt_653;   // oc8051_tb.v(104)
    output _cvpt_654;   // oc8051_tb.v(104)
    output _cvpt_655;   // oc8051_tb.v(104)
    output _cvpt_656;   // oc8051_tb.v(104)
    output _cvpt_657;   // oc8051_tb.v(104)
    output _cvpt_658;   // oc8051_tb.v(104)
    output _cvpt_659;   // oc8051_tb.v(104)
    output _cvpt_660;   // oc8051_tb.v(104)
    output _cvpt_661;   // oc8051_tb.v(104)
    output _cvpt_662;   // oc8051_tb.v(104)
    output _cvpt_663;   // oc8051_tb.v(104)
    output _cvpt_664;   // oc8051_tb.v(104)
    output _cvpt_665;   // oc8051_tb.v(104)
    output _cvpt_666;   // oc8051_tb.v(104)
    output _cvpt_667;   // oc8051_tb.v(104)
    output _cvpt_668;   // oc8051_tb.v(104)
    output _cvpt_669;   // oc8051_tb.v(104)
    output _cvpt_670;   // oc8051_tb.v(104)
    output _cvpt_671;   // oc8051_tb.v(104)
    output _cvpt_672;   // oc8051_tb.v(104)
    output _cvpt_673;   // oc8051_tb.v(104)
    output _cvpt_674;   // oc8051_tb.v(104)
    output _cvpt_675;   // oc8051_tb.v(104)
    output _cvpt_676;   // oc8051_tb.v(104)
    output _cvpt_677;   // oc8051_tb.v(104)
    output _cvpt_678;   // oc8051_tb.v(104)
    output _cvpt_679;   // oc8051_tb.v(104)
    output _cvpt_680;   // oc8051_tb.v(104)
    output _cvpt_681;   // oc8051_tb.v(104)
    output _cvpt_682;   // oc8051_tb.v(104)
    output _cvpt_683;   // oc8051_tb.v(104)
    output _cvpt_684;   // oc8051_tb.v(104)
    output _cvpt_685;   // oc8051_tb.v(104)
    output _cvpt_686;   // oc8051_tb.v(104)
    output _cvpt_687;   // oc8051_tb.v(104)
    output _cvpt_688;   // oc8051_tb.v(104)
    output _cvpt_689;   // oc8051_tb.v(104)
    output _cvpt_690;   // oc8051_tb.v(104)
    output _cvpt_691;   // oc8051_tb.v(104)
    output _cvpt_692;   // oc8051_tb.v(104)
    output _cvpt_693;   // oc8051_tb.v(104)
    output _cvpt_694;   // oc8051_tb.v(104)
    output _cvpt_695;   // oc8051_tb.v(104)
    output _cvpt_696;   // oc8051_tb.v(104)
    output _cvpt_697;   // oc8051_tb.v(104)
    output _cvpt_698;   // oc8051_tb.v(104)
    output _cvpt_699;   // oc8051_tb.v(104)
    output _cvpt_700;   // oc8051_tb.v(104)
    output _cvpt_701;   // oc8051_tb.v(104)
    output _cvpt_702;   // oc8051_tb.v(104)
    output _cvpt_703;   // oc8051_tb.v(104)
    output _cvpt_704;   // oc8051_tb.v(104)
    output _cvpt_705;   // oc8051_tb.v(104)
    output _cvpt_706;   // oc8051_tb.v(104)
    output _cvpt_707;   // oc8051_tb.v(104)
    output _cvpt_708;   // oc8051_tb.v(104)
    output _cvpt_709;   // oc8051_tb.v(104)
    output _cvpt_710;   // oc8051_tb.v(104)
    output _cvpt_711;   // oc8051_tb.v(104)
    output _cvpt_712;   // oc8051_tb.v(104)
    output _cvpt_713;   // oc8051_tb.v(104)
    output _cvpt_714;   // oc8051_tb.v(104)
    output _cvpt_715;   // oc8051_tb.v(104)
    output _cvpt_716;   // oc8051_tb.v(104)
    output _cvpt_717;   // oc8051_tb.v(104)
    output _cvpt_718;   // oc8051_tb.v(104)
    output _cvpt_719;   // oc8051_tb.v(104)
    output _cvpt_720;   // oc8051_tb.v(104)
    output _cvpt_721;   // oc8051_tb.v(104)
    output _cvpt_722;   // oc8051_tb.v(104)
    output _cvpt_723;   // oc8051_tb.v(104)
    output _cvpt_724;   // oc8051_tb.v(104)
    output _cvpt_725;   // oc8051_tb.v(104)
    output _cvpt_726;   // oc8051_tb.v(104)
    output _cvpt_727;   // oc8051_tb.v(104)
    output _cvpt_728;   // oc8051_tb.v(104)
    output _cvpt_729;   // oc8051_tb.v(104)
    output _cvpt_730;   // oc8051_tb.v(104)
    output _cvpt_731;   // oc8051_tb.v(104)
    output _cvpt_732;   // oc8051_tb.v(104)
    output _cvpt_733;   // oc8051_tb.v(104)
    output _cvpt_734;   // oc8051_tb.v(104)
    output _cvpt_735;   // oc8051_tb.v(104)
    output _cvpt_736;   // oc8051_tb.v(104)
    output _cvpt_737;   // oc8051_tb.v(104)
    output _cvpt_738;   // oc8051_tb.v(104)
    output _cvpt_739;   // oc8051_tb.v(104)
    output _cvpt_740;   // oc8051_tb.v(104)
    output _cvpt_741;   // oc8051_tb.v(104)
    output _cvpt_742;   // oc8051_tb.v(104)
    output _cvpt_743;   // oc8051_tb.v(104)
    output _cvpt_744;   // oc8051_tb.v(104)
    output _cvpt_745;   // oc8051_tb.v(104)
    output _cvpt_746;   // oc8051_tb.v(104)
    output _cvpt_747;   // oc8051_tb.v(104)
    output _cvpt_748;   // oc8051_tb.v(104)
    output _cvpt_749;   // oc8051_tb.v(104)
    output _cvpt_750;   // oc8051_tb.v(104)
    output _cvpt_751;   // oc8051_tb.v(104)
    output _cvpt_752;   // oc8051_tb.v(104)
    output _cvpt_753;   // oc8051_tb.v(104)
    output _cvpt_754;   // oc8051_tb.v(104)
    output _cvpt_755;   // oc8051_tb.v(104)
    output _cvpt_756;   // oc8051_tb.v(104)
    output _cvpt_757;   // oc8051_tb.v(104)
    output _cvpt_758;   // oc8051_tb.v(104)
    output _cvpt_759;   // oc8051_tb.v(104)
    output _cvpt_760;   // oc8051_tb.v(104)
    output _cvpt_761;   // oc8051_tb.v(104)
    output _cvpt_762;   // oc8051_tb.v(104)
    output _cvpt_763;   // oc8051_tb.v(104)
    output _cvpt_764;   // oc8051_tb.v(104)
    output _cvpt_765;   // oc8051_tb.v(104)
    output _cvpt_766;   // oc8051_tb.v(104)
    output _cvpt_767;   // oc8051_tb.v(104)
    output _cvpt_768;   // oc8051_tb.v(104)
    output _cvpt_769;   // oc8051_tb.v(104)
    output _cvpt_770;   // oc8051_tb.v(104)
    output _cvpt_771;   // oc8051_tb.v(104)
    output _cvpt_772;   // oc8051_tb.v(104)
    output _cvpt_773;   // oc8051_tb.v(104)
    output _cvpt_774;   // oc8051_tb.v(104)
    output _cvpt_775;   // oc8051_tb.v(104)
    output _cvpt_776;   // oc8051_tb.v(104)
    output _cvpt_777;   // oc8051_tb.v(104)
    output _cvpt_778;   // oc8051_tb.v(104)
    output _cvpt_779;   // oc8051_tb.v(104)
    output _cvpt_780;   // oc8051_tb.v(104)
    output _cvpt_781;   // oc8051_tb.v(104)
    output _cvpt_782;   // oc8051_tb.v(104)
    output _cvpt_783;   // oc8051_tb.v(104)
    output _cvpt_784;   // oc8051_tb.v(104)
    output _cvpt_785;   // oc8051_tb.v(104)
    output _cvpt_786;   // oc8051_tb.v(104)
    output _cvpt_787;   // oc8051_tb.v(104)
    output _cvpt_788;   // oc8051_tb.v(104)
    output _cvpt_789;   // oc8051_tb.v(104)
    output _cvpt_790;   // oc8051_tb.v(104)
    output _cvpt_791;   // oc8051_tb.v(104)
    output _cvpt_792;   // oc8051_tb.v(104)
    output _cvpt_793;   // oc8051_tb.v(104)
    output _cvpt_794;   // oc8051_tb.v(104)
    output _cvpt_795;   // oc8051_tb.v(104)
    output _cvpt_796;   // oc8051_tb.v(104)
    output _cvpt_797;   // oc8051_tb.v(104)
    output _cvpt_798;   // oc8051_tb.v(104)
    output _cvpt_799;   // oc8051_tb.v(104)
    output _cvpt_800;   // oc8051_tb.v(104)
    output _cvpt_801;   // oc8051_tb.v(104)
    output _cvpt_802;   // oc8051_tb.v(104)
    output _cvpt_803;   // oc8051_tb.v(104)
    output _cvpt_804;   // oc8051_tb.v(104)
    output _cvpt_805;   // oc8051_tb.v(104)
    output _cvpt_806;   // oc8051_tb.v(104)
    output _cvpt_807;   // oc8051_tb.v(104)
    output _cvpt_808;   // oc8051_tb.v(104)
    output _cvpt_809;   // oc8051_tb.v(104)
    output _cvpt_810;   // oc8051_tb.v(104)
    output _cvpt_811;   // oc8051_tb.v(104)
    output _cvpt_812;   // oc8051_tb.v(104)
    output _cvpt_813;   // oc8051_tb.v(104)
    output _cvpt_814;   // oc8051_tb.v(104)
    output _cvpt_815;   // oc8051_tb.v(104)
    output _cvpt_816;   // oc8051_tb.v(104)
    output _cvpt_817;   // oc8051_tb.v(104)
    output _cvpt_818;   // oc8051_tb.v(104)
    output _cvpt_819;   // oc8051_tb.v(104)
    output _cvpt_820;   // oc8051_tb.v(104)
    output _cvpt_821;   // oc8051_tb.v(104)
    output _cvpt_822;   // oc8051_tb.v(104)
    output _cvpt_823;   // oc8051_tb.v(104)
    output _cvpt_824;   // oc8051_tb.v(104)
    output _cvpt_825;   // oc8051_tb.v(104)
    output _cvpt_826;   // oc8051_tb.v(104)
    output _cvpt_827;   // oc8051_tb.v(104)
    output _cvpt_828;   // oc8051_tb.v(104)
    output _cvpt_829;   // oc8051_tb.v(104)
    output _cvpt_830;   // oc8051_tb.v(104)
    output _cvpt_831;   // oc8051_tb.v(104)
    output _cvpt_832;   // oc8051_tb.v(104)
    output _cvpt_833;   // oc8051_tb.v(104)
    output _cvpt_834;   // oc8051_tb.v(104)
    output _cvpt_835;   // oc8051_tb.v(104)
    output _cvpt_836;   // oc8051_tb.v(104)
    output _cvpt_837;   // oc8051_tb.v(104)
    output _cvpt_838;   // oc8051_tb.v(104)
    output _cvpt_839;   // oc8051_tb.v(104)
    output _cvpt_840;   // oc8051_tb.v(104)
    output _cvpt_841;   // oc8051_tb.v(104)
    output _cvpt_842;   // oc8051_tb.v(104)
    output _cvpt_843;   // oc8051_tb.v(104)
    output _cvpt_844;   // oc8051_tb.v(104)
    output _cvpt_845;   // oc8051_tb.v(104)
    output _cvpt_846;   // oc8051_tb.v(104)
    output _cvpt_847;   // oc8051_tb.v(104)
    output _cvpt_848;   // oc8051_tb.v(104)
    output _cvpt_849;   // oc8051_tb.v(104)
    output _cvpt_850;   // oc8051_tb.v(104)
    output _cvpt_851;   // oc8051_tb.v(104)
    output _cvpt_852;   // oc8051_tb.v(104)
    output _cvpt_853;   // oc8051_tb.v(104)
    output _cvpt_854;   // oc8051_tb.v(104)
    output _cvpt_855;   // oc8051_tb.v(104)
    output _cvpt_856;   // oc8051_tb.v(104)
    output _cvpt_857;   // oc8051_tb.v(104)
    output _cvpt_858;   // oc8051_tb.v(104)
    output _cvpt_859;   // oc8051_tb.v(104)
    output _cvpt_860;   // oc8051_tb.v(104)
    output _cvpt_861;   // oc8051_tb.v(104)
    output _cvpt_862;   // oc8051_tb.v(104)
    output _cvpt_863;   // oc8051_tb.v(104)
    output _cvpt_864;   // oc8051_tb.v(104)
    output _cvpt_865;   // oc8051_tb.v(104)
    output _cvpt_866;   // oc8051_tb.v(104)
    output _cvpt_867;   // oc8051_tb.v(104)
    output _cvpt_868;   // oc8051_tb.v(104)
    output _cvpt_869;   // oc8051_tb.v(104)
    output _cvpt_870;   // oc8051_tb.v(104)
    output _cvpt_871;   // oc8051_tb.v(104)
    output _cvpt_872;   // oc8051_tb.v(104)
    output _cvpt_873;   // oc8051_tb.v(104)
    output _cvpt_874;   // oc8051_tb.v(104)
    output _cvpt_875;   // oc8051_tb.v(104)
    output _cvpt_876;   // oc8051_tb.v(104)
    output _cvpt_877;   // oc8051_tb.v(104)
    output _cvpt_878;   // oc8051_tb.v(104)
    output _cvpt_879;   // oc8051_tb.v(104)
    output _cvpt_880;   // oc8051_tb.v(104)
    output _cvpt_881;   // oc8051_tb.v(104)
    output _cvpt_882;   // oc8051_tb.v(104)
    output _cvpt_883;   // oc8051_tb.v(104)
    output _cvpt_884;   // oc8051_tb.v(104)
    output _cvpt_885;   // oc8051_tb.v(104)
    output _cvpt_886;   // oc8051_tb.v(104)
    output _cvpt_887;   // oc8051_tb.v(104)
    output _cvpt_888;   // oc8051_tb.v(104)
    output _cvpt_889;   // oc8051_tb.v(104)
    output _cvpt_890;   // oc8051_tb.v(104)
    output _cvpt_891;   // oc8051_tb.v(104)
    output _cvpt_892;   // oc8051_tb.v(104)
    output _cvpt_893;   // oc8051_tb.v(104)
    output _cvpt_894;   // oc8051_tb.v(104)
    output _cvpt_895;   // oc8051_tb.v(104)
    output _cvpt_896;   // oc8051_tb.v(104)
    output _cvpt_897;   // oc8051_tb.v(104)
    output _cvpt_898;   // oc8051_tb.v(104)
    output _cvpt_899;   // oc8051_tb.v(104)
    output _cvpt_900;   // oc8051_tb.v(104)
    output _cvpt_901;   // oc8051_tb.v(104)
    output _cvpt_902;   // oc8051_tb.v(104)
    output _cvpt_903;   // oc8051_tb.v(104)
    output _cvpt_904;   // oc8051_tb.v(104)
    output _cvpt_905;   // oc8051_tb.v(104)
    output _cvpt_906;   // oc8051_tb.v(104)
    output _cvpt_907;   // oc8051_tb.v(104)
    output _cvpt_908;   // oc8051_tb.v(104)
    output _cvpt_909;   // oc8051_tb.v(104)
    output _cvpt_910;   // oc8051_tb.v(104)
    output _cvpt_911;   // oc8051_tb.v(104)
    output _cvpt_912;   // oc8051_tb.v(104)
    output _cvpt_913;   // oc8051_tb.v(104)
    output _cvpt_914;   // oc8051_tb.v(104)
    output _cvpt_915;   // oc8051_tb.v(104)
    output _cvpt_916;   // oc8051_tb.v(104)
    output _cvpt_917;   // oc8051_tb.v(104)
    output _cvpt_918;   // oc8051_tb.v(104)
    output _cvpt_919;   // oc8051_tb.v(104)
    output _cvpt_920;   // oc8051_tb.v(104)
    output _cvpt_921;   // oc8051_tb.v(104)
    output _cvpt_922;   // oc8051_tb.v(104)
    output _cvpt_923;   // oc8051_tb.v(104)
    output _cvpt_924;   // oc8051_tb.v(104)
    output _cvpt_925;   // oc8051_tb.v(104)
    output _cvpt_926;   // oc8051_tb.v(104)
    output _cvpt_927;   // oc8051_tb.v(104)
    output _cvpt_928;   // oc8051_tb.v(104)
    output _cvpt_929;   // oc8051_tb.v(104)
    output _cvpt_930;   // oc8051_tb.v(104)
    output _cvpt_931;   // oc8051_tb.v(104)
    output _cvpt_932;   // oc8051_tb.v(104)
    output _cvpt_933;   // oc8051_tb.v(104)
    output _cvpt_934;   // oc8051_tb.v(104)
    output _cvpt_935;   // oc8051_tb.v(104)
    output _cvpt_936;   // oc8051_tb.v(104)
    output _cvpt_937;   // oc8051_tb.v(104)
    output _cvpt_938;   // oc8051_tb.v(104)
    output _cvpt_939;   // oc8051_tb.v(104)
    output _cvpt_940;   // oc8051_tb.v(104)
    output _cvpt_941;   // oc8051_tb.v(104)
    output _cvpt_942;   // oc8051_tb.v(104)
    output _cvpt_943;   // oc8051_tb.v(104)
    output _cvpt_944;   // oc8051_tb.v(104)
    output _cvpt_945;   // oc8051_tb.v(104)
    output _cvpt_946;   // oc8051_tb.v(104)
    output _cvpt_947;   // oc8051_tb.v(104)
    output _cvpt_948;   // oc8051_tb.v(104)
    output _cvpt_949;   // oc8051_tb.v(104)
    output _cvpt_950;   // oc8051_tb.v(104)
    output _cvpt_951;   // oc8051_tb.v(104)
    output _cvpt_952;   // oc8051_tb.v(104)
    output _cvpt_953;   // oc8051_tb.v(104)
    output _cvpt_954;   // oc8051_tb.v(104)
    output _cvpt_955;   // oc8051_tb.v(104)
    output _cvpt_956;   // oc8051_tb.v(104)
    output _cvpt_957;   // oc8051_tb.v(104)
    output _cvpt_958;   // oc8051_tb.v(104)
    output _cvpt_959;   // oc8051_tb.v(104)
    output _cvpt_960;   // oc8051_tb.v(104)
    output _cvpt_961;   // oc8051_tb.v(104)
    output _cvpt_962;   // oc8051_tb.v(104)
    output _cvpt_963;   // oc8051_tb.v(104)
    output _cvpt_964;   // oc8051_tb.v(104)
    output _cvpt_965;   // oc8051_tb.v(104)
    output _cvpt_966;   // oc8051_tb.v(104)
    output _cvpt_967;   // oc8051_tb.v(104)
    output _cvpt_968;   // oc8051_tb.v(104)
    output _cvpt_969;   // oc8051_tb.v(104)
    output _cvpt_970;   // oc8051_tb.v(104)
    output _cvpt_971;   // oc8051_tb.v(104)
    output _cvpt_972;   // oc8051_tb.v(104)
    output _cvpt_973;   // oc8051_tb.v(104)
    output _cvpt_974;   // oc8051_tb.v(104)
    output _cvpt_975;   // oc8051_tb.v(104)
    output _cvpt_976;   // oc8051_tb.v(104)
    output _cvpt_977;   // oc8051_tb.v(104)
    output _cvpt_978;   // oc8051_tb.v(104)
    output _cvpt_979;   // oc8051_tb.v(104)
    output _cvpt_980;   // oc8051_tb.v(104)
    output _cvpt_981;   // oc8051_tb.v(104)
    output _cvpt_982;   // oc8051_tb.v(104)
    output _cvpt_983;   // oc8051_tb.v(104)
    output _cvpt_984;   // oc8051_tb.v(104)
    output _cvpt_985;   // oc8051_tb.v(104)
    output _cvpt_986;   // oc8051_tb.v(104)
    output _cvpt_987;   // oc8051_tb.v(104)
    output _cvpt_988;   // oc8051_tb.v(104)
    output _cvpt_989;   // oc8051_tb.v(104)
    output _cvpt_990;   // oc8051_tb.v(104)
    output _cvpt_991;   // oc8051_tb.v(104)
    output _cvpt_992;   // oc8051_tb.v(104)
    output _cvpt_993;   // oc8051_tb.v(104)
    output _cvpt_994;   // oc8051_tb.v(104)
    output _cvpt_995;   // oc8051_tb.v(104)
    output _cvpt_996;   // oc8051_tb.v(104)
    output _cvpt_997;   // oc8051_tb.v(104)
    output _cvpt_998;   // oc8051_tb.v(104)
    output _cvpt_999;   // oc8051_tb.v(104)
    output _cvpt_1000;   // oc8051_tb.v(104)
    output _cvpt_1001;   // oc8051_tb.v(104)
    output _cvpt_1002;   // oc8051_tb.v(104)
    output _cvpt_1003;   // oc8051_tb.v(104)
    output _cvpt_1004;   // oc8051_tb.v(104)
    output _cvpt_1005;   // oc8051_tb.v(104)
    output _cvpt_1006;   // oc8051_tb.v(104)
    output _cvpt_1007;   // oc8051_tb.v(104)
    output _cvpt_1008;   // oc8051_tb.v(104)
    output _cvpt_1009;   // oc8051_tb.v(104)
    output _cvpt_1010;   // oc8051_tb.v(104)
    output _cvpt_1011;   // oc8051_tb.v(104)
    output _cvpt_1012;   // oc8051_tb.v(104)
    output _cvpt_1013;   // oc8051_tb.v(104)
    output _cvpt_1014;   // oc8051_tb.v(104)
    output _cvpt_1015;   // oc8051_tb.v(104)
    output _cvpt_1016;   // oc8051_tb.v(104)
    output _cvpt_1017;   // oc8051_tb.v(104)
    output _cvpt_1018;   // oc8051_tb.v(104)
    output _cvpt_1019;   // oc8051_tb.v(104)
    output _cvpt_1020;   // oc8051_tb.v(104)
    output _cvpt_1021;   // oc8051_tb.v(104)
    output _cvpt_1022;   // oc8051_tb.v(104)
    output _cvpt_1023;   // oc8051_tb.v(104)
    output _cvpt_1024;   // oc8051_tb.v(104)
    output _cvpt_1025;   // oc8051_tb.v(104)
    output _cvpt_1026;   // oc8051_tb.v(104)
    output _cvpt_1027;   // oc8051_tb.v(104)
    output _cvpt_1028;   // oc8051_tb.v(104)
    output _cvpt_1029;   // oc8051_tb.v(104)
    output _cvpt_1030;   // oc8051_tb.v(104)
    output _cvpt_1031;   // oc8051_tb.v(104)
    output _cvpt_1032;   // oc8051_tb.v(104)
    output _cvpt_1033;   // oc8051_tb.v(104)
    output _cvpt_1034;   // oc8051_tb.v(104)
    output _cvpt_1035;   // oc8051_tb.v(104)
    output _cvpt_1036;   // oc8051_tb.v(104)
    output _cvpt_1037;   // oc8051_tb.v(104)
    output _cvpt_1038;   // oc8051_tb.v(104)
    output _cvpt_1039;   // oc8051_tb.v(104)
    output _cvpt_1040;   // oc8051_tb.v(104)
    output _cvpt_1041;   // oc8051_tb.v(104)
    output _cvpt_1042;   // oc8051_tb.v(104)
    output _cvpt_1043;   // oc8051_tb.v(104)
    output _cvpt_1044;   // oc8051_tb.v(104)
    output _cvpt_1045;   // oc8051_tb.v(104)
    output _cvpt_1046;   // oc8051_tb.v(104)
    output _cvpt_1047;   // oc8051_tb.v(104)
    output _cvpt_1048;   // oc8051_tb.v(104)
    output _cvpt_1049;   // oc8051_tb.v(104)
    output _cvpt_1050;   // oc8051_tb.v(104)
    output _cvpt_1051;   // oc8051_tb.v(104)
    output _cvpt_1052;   // oc8051_tb.v(104)
    output _cvpt_1053;   // oc8051_tb.v(104)
    output _cvpt_1054;   // oc8051_tb.v(104)
    output _cvpt_1055;   // oc8051_tb.v(104)
    output _cvpt_1056;   // oc8051_tb.v(104)
    output _cvpt_1057;   // oc8051_tb.v(104)
    output _cvpt_1058;   // oc8051_tb.v(104)
    output _cvpt_1059;   // oc8051_tb.v(104)
    output _cvpt_1060;   // oc8051_tb.v(104)
    output _cvpt_1061;   // oc8051_tb.v(104)
    output _cvpt_1062;   // oc8051_tb.v(104)
    output _cvpt_1063;   // oc8051_tb.v(104)
    output _cvpt_1064;   // oc8051_tb.v(104)
    output _cvpt_1065;   // oc8051_tb.v(104)
    output _cvpt_1066;   // oc8051_tb.v(104)
    output _cvpt_1067;   // oc8051_tb.v(104)
    output _cvpt_1068;   // oc8051_tb.v(104)
    output _cvpt_1069;   // oc8051_tb.v(104)
    output _cvpt_1070;   // oc8051_tb.v(104)
    output _cvpt_1071;   // oc8051_tb.v(104)
    output _cvpt_1072;   // oc8051_tb.v(104)
    output _cvpt_1073;   // oc8051_tb.v(104)
    output _cvpt_1074;   // oc8051_tb.v(104)
    output _cvpt_1075;   // oc8051_tb.v(104)
    output _cvpt_1076;   // oc8051_tb.v(104)
    output _cvpt_1077;   // oc8051_tb.v(104)
    output _cvpt_1078;   // oc8051_tb.v(104)
    output _cvpt_1079;   // oc8051_tb.v(104)
    output _cvpt_1080;   // oc8051_tb.v(104)
    output _cvpt_1081;   // oc8051_tb.v(104)
    output _cvpt_1082;   // oc8051_tb.v(104)
    output _cvpt_1083;   // oc8051_tb.v(104)
    output _cvpt_1084;   // oc8051_tb.v(104)
    output _cvpt_1085;   // oc8051_tb.v(104)
    output _cvpt_1086;   // oc8051_tb.v(104)
    output _cvpt_1087;   // oc8051_tb.v(104)
    output _cvpt_1088;   // oc8051_tb.v(104)
    output _cvpt_1089;   // oc8051_tb.v(104)
    output _cvpt_1090;   // oc8051_tb.v(104)
    output _cvpt_1091;   // oc8051_tb.v(104)
    output _cvpt_1092;   // oc8051_tb.v(104)
    output _cvpt_1093;   // oc8051_tb.v(104)
    output _cvpt_1094;   // oc8051_tb.v(104)
    output _cvpt_1095;   // oc8051_tb.v(104)
    output _cvpt_1096;   // oc8051_tb.v(104)
    output _cvpt_1097;   // oc8051_tb.v(104)
    output _cvpt_1098;   // oc8051_tb.v(104)
    output _cvpt_1099;   // oc8051_tb.v(104)
    output _cvpt_1100;   // oc8051_tb.v(104)
    output _cvpt_1101;   // oc8051_tb.v(104)
    output _cvpt_1102;   // oc8051_tb.v(104)
    output _cvpt_1103;   // oc8051_tb.v(104)
    output _cvpt_1104;   // oc8051_tb.v(104)
    output _cvpt_1105;   // oc8051_tb.v(104)
    output _cvpt_1106;   // oc8051_tb.v(104)
    output _cvpt_1107;   // oc8051_tb.v(104)
    output _cvpt_1108;   // oc8051_tb.v(104)
    output _cvpt_1109;   // oc8051_tb.v(104)
    output _cvpt_1110;   // oc8051_tb.v(104)
    output _cvpt_1111;   // oc8051_tb.v(104)
    output _cvpt_1112;   // oc8051_tb.v(104)
    output _cvpt_1113;   // oc8051_tb.v(104)
    output _cvpt_1114;   // oc8051_tb.v(104)
    output _cvpt_1115;   // oc8051_tb.v(104)
    output _cvpt_1116;   // oc8051_tb.v(104)
    output _cvpt_1117;   // oc8051_tb.v(104)
    output _cvpt_1118;   // oc8051_tb.v(104)
    output _cvpt_1119;   // oc8051_tb.v(104)
    output _cvpt_1120;   // oc8051_tb.v(104)
    output _cvpt_1121;   // oc8051_tb.v(104)
    output _cvpt_1122;   // oc8051_tb.v(104)
    output _cvpt_1123;   // oc8051_tb.v(104)
    output _cvpt_1124;   // oc8051_tb.v(104)
    output _cvpt_1125;   // oc8051_tb.v(104)
    output _cvpt_1126;   // oc8051_tb.v(104)
    output _cvpt_1127;   // oc8051_tb.v(104)
    output _cvpt_1128;   // oc8051_tb.v(104)
    output _cvpt_1129;   // oc8051_tb.v(104)
    output _cvpt_1130;   // oc8051_tb.v(104)
    output _cvpt_1131;   // oc8051_tb.v(104)
    output _cvpt_1132;   // oc8051_tb.v(104)
    output _cvpt_1133;   // oc8051_tb.v(104)
    output _cvpt_1134;   // oc8051_tb.v(104)
    output _cvpt_1135;   // oc8051_tb.v(104)
    output _cvpt_1136;   // oc8051_tb.v(104)
    output _cvpt_1137;   // oc8051_tb.v(104)
    output _cvpt_1138;   // oc8051_tb.v(104)
    output _cvpt_1139;   // oc8051_tb.v(104)
    output _cvpt_1140;   // oc8051_tb.v(104)
    output _cvpt_1141;   // oc8051_tb.v(104)
    output _cvpt_1142;   // oc8051_tb.v(104)
    output _cvpt_1143;   // oc8051_tb.v(104)
    output _cvpt_1144;   // oc8051_tb.v(104)
    output _cvpt_1145;   // oc8051_tb.v(104)
    output _cvpt_1146;   // oc8051_tb.v(104)
    output _cvpt_1147;   // oc8051_tb.v(104)
    output _cvpt_1148;   // oc8051_tb.v(104)
    output _cvpt_1149;   // oc8051_tb.v(104)
    output _cvpt_1150;   // oc8051_tb.v(104)
    output _cvpt_1151;   // oc8051_tb.v(104)
    output _cvpt_1152;   // oc8051_tb.v(104)
    output _cvpt_1153;   // oc8051_tb.v(104)
    output _cvpt_1154;   // oc8051_tb.v(104)
    output _cvpt_1155;   // oc8051_tb.v(104)
    output _cvpt_1156;   // oc8051_tb.v(104)
    output _cvpt_1157;   // oc8051_tb.v(104)
    output _cvpt_1158;   // oc8051_tb.v(104)
    output _cvpt_1159;   // oc8051_tb.v(104)
    output _cvpt_1160;   // oc8051_tb.v(104)
    output _cvpt_1161;   // oc8051_tb.v(104)
    output _cvpt_1162;   // oc8051_tb.v(104)
    output _cvpt_1163;   // oc8051_tb.v(104)
    output _cvpt_1164;   // oc8051_tb.v(104)
    output _cvpt_1165;   // oc8051_tb.v(104)
    output _cvpt_1166;   // oc8051_tb.v(104)
    output _cvpt_1167;   // oc8051_tb.v(104)
    output _cvpt_1168;   // oc8051_tb.v(104)
    output _cvpt_1169;   // oc8051_tb.v(104)
    output _cvpt_1170;   // oc8051_tb.v(104)
    output _cvpt_1171;   // oc8051_tb.v(104)
    output _cvpt_1172;   // oc8051_tb.v(104)
    output _cvpt_1173;   // oc8051_tb.v(104)
    output _cvpt_1174;   // oc8051_tb.v(104)
    output _cvpt_1175;   // oc8051_tb.v(104)
    output _cvpt_1176;   // oc8051_tb.v(104)
    output _cvpt_1177;   // oc8051_tb.v(104)
    output _cvpt_1178;   // oc8051_tb.v(104)
    output _cvpt_1179;   // oc8051_tb.v(104)
    output _cvpt_1180;   // oc8051_tb.v(104)
    output _cvpt_1181;   // oc8051_tb.v(104)
    output _cvpt_1182;   // oc8051_tb.v(104)
    output _cvpt_1183;   // oc8051_tb.v(104)
    output _cvpt_1184;   // oc8051_tb.v(104)
    output _cvpt_1185;   // oc8051_tb.v(104)
    output _cvpt_1186;   // oc8051_tb.v(104)
    output _cvpt_1187;   // oc8051_tb.v(104)
    output _cvpt_1188;   // oc8051_tb.v(104)
    output _cvpt_1189;   // oc8051_tb.v(104)
    output _cvpt_1190;   // oc8051_tb.v(104)
    output _cvpt_1191;   // oc8051_tb.v(104)
    output _cvpt_1192;   // oc8051_tb.v(104)
    output _cvpt_1193;   // oc8051_tb.v(104)
    output _cvpt_1194;   // oc8051_tb.v(104)
    output _cvpt_1195;   // oc8051_tb.v(104)
    output _cvpt_1196;   // oc8051_tb.v(104)
    output _cvpt_1197;   // oc8051_tb.v(104)
    output _cvpt_1198;   // oc8051_tb.v(104)
    output _cvpt_1199;   // oc8051_tb.v(104)
    output _cvpt_1200;   // oc8051_tb.v(104)
    output _cvpt_1201;   // oc8051_tb.v(104)
    output _cvpt_1202;   // oc8051_tb.v(104)
    output _cvpt_1203;   // oc8051_tb.v(104)
    output _cvpt_1204;   // oc8051_tb.v(104)
    output _cvpt_1205;   // oc8051_tb.v(104)
    output _cvpt_1206;   // oc8051_tb.v(104)
    output _cvpt_1207;   // oc8051_tb.v(104)
    output _cvpt_1208;   // oc8051_tb.v(104)
    output _cvpt_1209;   // oc8051_tb.v(104)
    output _cvpt_1210;   // oc8051_tb.v(104)
    output _cvpt_1211;   // oc8051_tb.v(104)
    output _cvpt_1212;   // oc8051_tb.v(104)
    output _cvpt_1213;   // oc8051_tb.v(104)
    output _cvpt_1214;   // oc8051_tb.v(104)
    output _cvpt_1215;   // oc8051_tb.v(104)
    output _cvpt_1216;   // oc8051_tb.v(104)
    output _cvpt_1217;   // oc8051_tb.v(104)
    output _cvpt_1218;   // oc8051_tb.v(104)
    output _cvpt_1219;   // oc8051_tb.v(104)
    output _cvpt_1220;   // oc8051_tb.v(104)
    output _cvpt_1221;   // oc8051_tb.v(104)
    output _cvpt_1222;   // oc8051_tb.v(104)
    output _cvpt_1223;   // oc8051_tb.v(104)
    output _cvpt_1224;   // oc8051_tb.v(104)
    output _cvpt_1225;   // oc8051_tb.v(104)
    output _cvpt_1226;   // oc8051_tb.v(104)
    output _cvpt_1227;   // oc8051_tb.v(104)
    output _cvpt_1228;   // oc8051_tb.v(104)
    output _cvpt_1229;   // oc8051_tb.v(104)
    output _cvpt_1230;   // oc8051_tb.v(104)
    output _cvpt_1231;   // oc8051_tb.v(104)
    output _cvpt_1232;   // oc8051_tb.v(104)
    output _cvpt_1233;   // oc8051_tb.v(104)
    output _cvpt_1234;   // oc8051_tb.v(104)
    output _cvpt_1235;   // oc8051_tb.v(104)
    output _cvpt_1236;   // oc8051_tb.v(104)
    output _cvpt_1237;   // oc8051_tb.v(104)
    output _cvpt_1238;   // oc8051_tb.v(104)
    output _cvpt_1239;   // oc8051_tb.v(104)
    output _cvpt_1240;   // oc8051_tb.v(104)
    output _cvpt_1241;   // oc8051_tb.v(104)
    output _cvpt_1242;   // oc8051_tb.v(104)
    output _cvpt_1243;   // oc8051_tb.v(104)
    output _cvpt_1244;   // oc8051_tb.v(104)
    output _cvpt_1245;   // oc8051_tb.v(104)
    output _cvpt_1246;   // oc8051_tb.v(104)
    output _cvpt_1247;   // oc8051_tb.v(104)
    output _cvpt_1248;   // oc8051_tb.v(104)
    output _cvpt_1249;   // oc8051_tb.v(104)
    output _cvpt_1250;   // oc8051_tb.v(104)
    output _cvpt_1251;   // oc8051_tb.v(104)
    output _cvpt_1252;   // oc8051_tb.v(104)
    output _cvpt_1253;   // oc8051_tb.v(104)
    output _cvpt_1254;   // oc8051_tb.v(104)
    output _cvpt_1255;   // oc8051_tb.v(104)
    output _cvpt_1256;   // oc8051_tb.v(104)
    output _cvpt_1257;   // oc8051_tb.v(104)
    output _cvpt_1258;   // oc8051_tb.v(104)
    output _cvpt_1259;   // oc8051_tb.v(104)
    output _cvpt_1260;   // oc8051_tb.v(104)
    output _cvpt_1261;   // oc8051_tb.v(104)
    output _cvpt_1262;   // oc8051_tb.v(104)
    output _cvpt_1263;   // oc8051_tb.v(104)
    output _cvpt_1264;   // oc8051_tb.v(104)
    output _cvpt_1265;   // oc8051_tb.v(104)
    output _cvpt_1266;   // oc8051_tb.v(104)
    output _cvpt_1267;   // oc8051_tb.v(104)
    output _cvpt_1268;   // oc8051_tb.v(104)
    output _cvpt_1269;   // oc8051_tb.v(104)
    output _cvpt_1270;   // oc8051_tb.v(104)
    output _cvpt_1271;   // oc8051_tb.v(104)
    output _cvpt_1272;   // oc8051_tb.v(104)
    output _cvpt_1273;   // oc8051_tb.v(104)
    output _cvpt_1274;   // oc8051_tb.v(104)
    output _cvpt_1275;   // oc8051_tb.v(104)
    output _cvpt_1276;   // oc8051_tb.v(104)
    output _cvpt_1277;   // oc8051_tb.v(104)
    output _cvpt_1278;   // oc8051_tb.v(104)
    output _cvpt_1279;   // oc8051_tb.v(104)
    output _cvpt_1280;   // oc8051_tb.v(104)
    output _cvpt_1281;   // oc8051_tb.v(104)
    output _cvpt_1282;   // oc8051_tb.v(104)
    output _cvpt_1283;   // oc8051_tb.v(104)
    output _cvpt_1284;   // oc8051_tb.v(104)
    output _cvpt_1285;   // oc8051_tb.v(104)
    output _cvpt_1286;   // oc8051_tb.v(104)
    output _cvpt_1287;   // oc8051_tb.v(104)
    output _cvpt_1288;   // oc8051_tb.v(104)
    output _cvpt_1289;   // oc8051_tb.v(104)
    output _cvpt_1290;   // oc8051_tb.v(104)
    output _cvpt_1291;   // oc8051_tb.v(104)
    output _cvpt_1292;   // oc8051_tb.v(104)
    output _cvpt_1293;   // oc8051_tb.v(104)
    output _cvpt_1294;   // oc8051_tb.v(104)
    output _cvpt_1295;   // oc8051_tb.v(104)
    output _cvpt_1296;   // oc8051_tb.v(104)
    output _cvpt_1297;   // oc8051_tb.v(104)
    output _cvpt_1298;   // oc8051_tb.v(104)
    output _cvpt_1299;   // oc8051_tb.v(104)
    output _cvpt_1300;   // oc8051_tb.v(104)
    output _cvpt_1301;   // oc8051_tb.v(104)
    output _cvpt_1302;   // oc8051_tb.v(104)
    output _cvpt_1303;   // oc8051_tb.v(104)
    output _cvpt_1304;   // oc8051_tb.v(104)
    output _cvpt_1305;   // oc8051_tb.v(104)
    output _cvpt_1306;   // oc8051_tb.v(104)
    output _cvpt_1307;   // oc8051_tb.v(104)
    output _cvpt_1308;   // oc8051_tb.v(104)
    output _cvpt_1309;   // oc8051_tb.v(104)
    output _cvpt_1310;   // oc8051_tb.v(104)
    output _cvpt_1311;   // oc8051_tb.v(104)
    output _cvpt_1312;   // oc8051_tb.v(104)
    output _cvpt_1313;   // oc8051_tb.v(104)
    output _cvpt_1314;   // oc8051_tb.v(104)
    output _cvpt_1315;   // oc8051_tb.v(104)
    output _cvpt_1316;   // oc8051_tb.v(104)
    output _cvpt_1317;   // oc8051_tb.v(104)
    output _cvpt_1318;   // oc8051_tb.v(104)
    output _cvpt_1319;   // oc8051_tb.v(104)
    output _cvpt_1320;   // oc8051_tb.v(104)
    output _cvpt_1321;   // oc8051_tb.v(104)
    output _cvpt_1322;   // oc8051_tb.v(104)
    output _cvpt_1323;   // oc8051_tb.v(104)
    output _cvpt_1324;   // oc8051_tb.v(104)
    output _cvpt_1325;   // oc8051_tb.v(104)
    output _cvpt_1326;   // oc8051_tb.v(104)
    output _cvpt_1327;   // oc8051_tb.v(104)
    output _cvpt_1328;   // oc8051_tb.v(104)
    output _cvpt_1329;   // oc8051_tb.v(104)
    output _cvpt_1330;   // oc8051_tb.v(104)
    output _cvpt_1331;   // oc8051_tb.v(104)
    output _cvpt_1332;   // oc8051_tb.v(104)
    output _cvpt_1333;   // oc8051_tb.v(104)
    output _cvpt_1334;   // oc8051_tb.v(104)
    output _cvpt_1335;   // oc8051_tb.v(104)
    output _cvpt_1336;   // oc8051_tb.v(104)
    output _cvpt_1337;   // oc8051_tb.v(104)
    output _cvpt_1338;   // oc8051_tb.v(104)
    output _cvpt_1339;   // oc8051_tb.v(104)
    output _cvpt_1340;   // oc8051_tb.v(104)
    output _cvpt_1341;   // oc8051_tb.v(104)
    output _cvpt_1342;   // oc8051_tb.v(104)
    output _cvpt_1343;   // oc8051_tb.v(104)
    output _cvpt_1344;   // oc8051_tb.v(104)
    output _cvpt_1345;   // oc8051_tb.v(104)
    output _cvpt_1346;   // oc8051_tb.v(104)
    output _cvpt_1347;   // oc8051_tb.v(104)
    output _cvpt_1348;   // oc8051_tb.v(104)
    output _cvpt_1349;   // oc8051_tb.v(104)
    output _cvpt_1350;   // oc8051_tb.v(104)
    output _cvpt_1351;   // oc8051_tb.v(104)
    output _cvpt_1352;   // oc8051_tb.v(104)
    output _cvpt_1353;   // oc8051_tb.v(104)
    output _cvpt_1354;   // oc8051_tb.v(104)
    output _cvpt_1355;   // oc8051_tb.v(104)
    output _cvpt_1356;   // oc8051_tb.v(104)
    output _cvpt_1357;   // oc8051_tb.v(104)
    output _cvpt_1358;   // oc8051_tb.v(104)
    output _cvpt_1359;   // oc8051_tb.v(104)
    output _cvpt_1360;   // oc8051_tb.v(104)
    output _cvpt_1361;   // oc8051_tb.v(104)
    output _cvpt_1362;   // oc8051_tb.v(104)
    output _cvpt_1363;   // oc8051_tb.v(104)
    output _cvpt_1364;   // oc8051_tb.v(104)
    output _cvpt_1365;   // oc8051_tb.v(104)
    output _cvpt_1366;   // oc8051_tb.v(104)
    output _cvpt_1367;   // oc8051_tb.v(104)
    output _cvpt_1368;   // oc8051_tb.v(104)
    output _cvpt_1369;   // oc8051_tb.v(104)
    output _cvpt_1370;   // oc8051_tb.v(104)
    output _cvpt_1371;   // oc8051_tb.v(104)
    output _cvpt_1372;   // oc8051_tb.v(104)
    output _cvpt_1373;   // oc8051_tb.v(104)
    output _cvpt_1374;   // oc8051_tb.v(104)
    output _cvpt_1375;   // oc8051_tb.v(104)
    output _cvpt_1376;   // oc8051_tb.v(104)
    output _cvpt_1377;   // oc8051_tb.v(104)
    output _cvpt_1378;   // oc8051_tb.v(104)
    output _cvpt_1379;   // oc8051_tb.v(104)
    output _cvpt_1380;   // oc8051_tb.v(104)
    output _cvpt_1381;   // oc8051_tb.v(104)
    output _cvpt_1382;   // oc8051_tb.v(104)
    output _cvpt_1383;   // oc8051_tb.v(104)
    output _cvpt_1384;   // oc8051_tb.v(104)
    output _cvpt_1385;   // oc8051_tb.v(104)
    output _cvpt_1386;   // oc8051_tb.v(104)
    output _cvpt_1387;   // oc8051_tb.v(104)
    output _cvpt_1388;   // oc8051_tb.v(104)
    output _cvpt_1389;   // oc8051_tb.v(104)
    output _cvpt_1390;   // oc8051_tb.v(104)
    output _cvpt_1391;   // oc8051_tb.v(104)
    output _cvpt_1392;   // oc8051_tb.v(104)
    output _cvpt_1393;   // oc8051_tb.v(104)
    output _cvpt_1394;   // oc8051_tb.v(104)
    output _cvpt_1395;   // oc8051_tb.v(104)
    output _cvpt_1396;   // oc8051_tb.v(104)
    output _cvpt_1397;   // oc8051_tb.v(104)
    output _cvpt_1398;   // oc8051_tb.v(104)
    output _cvpt_1399;   // oc8051_tb.v(104)
    output _cvpt_1400;   // oc8051_tb.v(104)
    output _cvpt_1401;   // oc8051_tb.v(104)
    output _cvpt_1402;   // oc8051_tb.v(104)
    output _cvpt_1403;   // oc8051_tb.v(104)
    output _cvpt_1404;   // oc8051_tb.v(104)
    output _cvpt_1405;   // oc8051_tb.v(104)
    output _cvpt_1406;   // oc8051_tb.v(104)
    output _cvpt_1407;   // oc8051_tb.v(104)
    output _cvpt_1408;   // oc8051_tb.v(104)
    output _cvpt_1409;   // oc8051_tb.v(104)
    output _cvpt_1410;   // oc8051_tb.v(104)
    output _cvpt_1411;   // oc8051_tb.v(104)
    output _cvpt_1412;   // oc8051_tb.v(104)
    output _cvpt_1413;   // oc8051_tb.v(104)
    output _cvpt_1414;   // oc8051_tb.v(104)
    output _cvpt_1415;   // oc8051_tb.v(104)
    output _cvpt_1416;   // oc8051_tb.v(104)
    output _cvpt_1417;   // oc8051_tb.v(104)
    output _cvpt_1418;   // oc8051_tb.v(104)
    output _cvpt_1419;   // oc8051_tb.v(104)
    output _cvpt_1420;   // oc8051_tb.v(104)
    output _cvpt_1421;   // oc8051_tb.v(104)
    output _cvpt_1422;   // oc8051_tb.v(104)
    output _cvpt_1423;   // oc8051_tb.v(104)
    output _cvpt_1424;   // oc8051_tb.v(104)
    output _cvpt_1425;   // oc8051_tb.v(104)
    output _cvpt_1426;   // oc8051_tb.v(104)
    output _cvpt_1427;   // oc8051_tb.v(104)
    output _cvpt_1428;   // oc8051_tb.v(104)
    output _cvpt_1429;   // oc8051_tb.v(104)
    output _cvpt_1430;   // oc8051_tb.v(104)
    output _cvpt_1431;   // oc8051_tb.v(104)
    output _cvpt_1432;   // oc8051_tb.v(104)
    output _cvpt_1433;   // oc8051_tb.v(104)
    output _cvpt_1434;   // oc8051_tb.v(104)
    output _cvpt_1435;   // oc8051_tb.v(104)
    output _cvpt_1436;   // oc8051_tb.v(104)
    output _cvpt_1437;   // oc8051_tb.v(104)
    output _cvpt_1438;   // oc8051_tb.v(104)
    output _cvpt_1439;   // oc8051_tb.v(104)
    output _cvpt_1440;   // oc8051_tb.v(104)
    output _cvpt_1441;   // oc8051_tb.v(104)
    output _cvpt_1442;   // oc8051_tb.v(104)
    output _cvpt_1443;   // oc8051_tb.v(104)
    output _cvpt_1444;   // oc8051_tb.v(104)
    output _cvpt_1445;   // oc8051_tb.v(104)
    output _cvpt_1446;   // oc8051_tb.v(104)
    output _cvpt_1447;   // oc8051_tb.v(104)
    output _cvpt_1448;   // oc8051_tb.v(104)
    output _cvpt_1449;   // oc8051_tb.v(104)
    output _cvpt_1450;   // oc8051_tb.v(104)
    output _cvpt_1451;   // oc8051_tb.v(104)
    output _cvpt_1452;   // oc8051_tb.v(104)
    output _cvpt_1453;   // oc8051_tb.v(104)
    output _cvpt_1454;   // oc8051_tb.v(104)
    output _cvpt_1455;   // oc8051_tb.v(104)
    output _cvpt_1456;   // oc8051_tb.v(104)
    output _cvpt_1457;   // oc8051_tb.v(104)
    output _cvpt_1458;   // oc8051_tb.v(104)
    output _cvpt_1459;   // oc8051_tb.v(104)
    output _cvpt_1460;   // oc8051_tb.v(104)
    output _cvpt_1461;   // oc8051_tb.v(104)
    output _cvpt_1462;   // oc8051_tb.v(104)
    output _cvpt_1463;   // oc8051_tb.v(104)
    output _cvpt_1464;   // oc8051_tb.v(104)
    output _cvpt_1465;   // oc8051_tb.v(104)
    output _cvpt_1466;   // oc8051_tb.v(104)
    output _cvpt_1467;   // oc8051_tb.v(104)
    output _cvpt_1468;   // oc8051_tb.v(104)
    output _cvpt_1469;   // oc8051_tb.v(104)
    output _cvpt_1470;   // oc8051_tb.v(104)
    output _cvpt_1471;   // oc8051_tb.v(104)
    output _cvpt_1472;   // oc8051_tb.v(104)
    output _cvpt_1473;   // oc8051_tb.v(104)
    output _cvpt_1474;   // oc8051_tb.v(104)
    output _cvpt_1475;   // oc8051_tb.v(104)
    output _cvpt_1476;   // oc8051_tb.v(104)
    output _cvpt_1477;   // oc8051_tb.v(104)
    output _cvpt_1478;   // oc8051_tb.v(104)
    output _cvpt_1479;   // oc8051_tb.v(104)
    output _cvpt_1480;   // oc8051_tb.v(104)
    output _cvpt_1481;   // oc8051_tb.v(104)
    output _cvpt_1482;   // oc8051_tb.v(104)
    output _cvpt_1483;   // oc8051_tb.v(104)
    output _cvpt_1484;   // oc8051_tb.v(104)
    output _cvpt_1485;   // oc8051_tb.v(104)
    output _cvpt_1486;   // oc8051_tb.v(104)
    output _cvpt_1487;   // oc8051_tb.v(104)
    output _cvpt_1488;   // oc8051_tb.v(104)
    output _cvpt_1489;   // oc8051_tb.v(104)
    output _cvpt_1490;   // oc8051_tb.v(104)
    output _cvpt_1491;   // oc8051_tb.v(104)
    output _cvpt_1492;   // oc8051_tb.v(104)
    output _cvpt_1493;   // oc8051_tb.v(104)
    output _cvpt_1494;   // oc8051_tb.v(104)
    output _cvpt_1495;   // oc8051_tb.v(104)
    output _cvpt_1496;   // oc8051_tb.v(104)
    output _cvpt_1497;   // oc8051_tb.v(104)
    output _cvpt_1498;   // oc8051_tb.v(104)
    output _cvpt_1499;   // oc8051_tb.v(104)
    output _cvpt_1500;   // oc8051_tb.v(104)
    output _cvpt_1501;   // oc8051_tb.v(104)
    output _cvpt_1502;   // oc8051_tb.v(104)
    output _cvpt_1503;   // oc8051_tb.v(104)
    output _cvpt_1504;   // oc8051_tb.v(104)
    output _cvpt_1505;   // oc8051_tb.v(104)
    output _cvpt_1506;   // oc8051_tb.v(104)
    output _cvpt_1507;   // oc8051_tb.v(104)
    output _cvpt_1508;   // oc8051_tb.v(104)
    output _cvpt_1509;   // oc8051_tb.v(104)
    output _cvpt_1510;   // oc8051_tb.v(104)
    output _cvpt_1511;   // oc8051_tb.v(104)
    output _cvpt_1512;   // oc8051_tb.v(104)
    output _cvpt_1513;   // oc8051_tb.v(104)
    output _cvpt_1514;   // oc8051_tb.v(104)
    output _cvpt_1515;   // oc8051_tb.v(104)
    output _cvpt_1516;   // oc8051_tb.v(104)
    output _cvpt_1517;   // oc8051_tb.v(104)
    output _cvpt_1518;   // oc8051_tb.v(104)
    output _cvpt_1519;   // oc8051_tb.v(104)
    output _cvpt_1520;   // oc8051_tb.v(104)
    output _cvpt_1521;   // oc8051_tb.v(104)
    output _cvpt_1522;   // oc8051_tb.v(104)
    output _cvpt_1523;   // oc8051_tb.v(104)
    output _cvpt_1524;   // oc8051_tb.v(104)
    output _cvpt_1525;   // oc8051_tb.v(104)
    output _cvpt_1526;   // oc8051_tb.v(104)
    output _cvpt_1527;   // oc8051_tb.v(104)
    output _cvpt_1528;   // oc8051_tb.v(104)
    output _cvpt_1529;   // oc8051_tb.v(104)
    output _cvpt_1530;   // oc8051_tb.v(104)
    output _cvpt_1531;   // oc8051_tb.v(104)
    output _cvpt_1532;   // oc8051_tb.v(104)
    output _cvpt_1533;   // oc8051_tb.v(104)
    output _cvpt_1534;   // oc8051_tb.v(104)
    output _cvpt_1535;   // oc8051_tb.v(104)
    output _cvpt_1536;   // oc8051_tb.v(104)
    output _cvpt_1537;   // oc8051_tb.v(104)
    output _cvpt_1538;   // oc8051_tb.v(104)
    output _cvpt_1539;   // oc8051_tb.v(104)
    output _cvpt_1540;   // oc8051_tb.v(104)
    output _cvpt_1541;   // oc8051_tb.v(104)
    output _cvpt_1542;   // oc8051_tb.v(104)
    output _cvpt_1543;   // oc8051_tb.v(104)
    output _cvpt_1544;   // oc8051_tb.v(104)
    output _cvpt_1545;   // oc8051_tb.v(104)
    output _cvpt_1546;   // oc8051_tb.v(104)
    output _cvpt_1547;   // oc8051_tb.v(104)
    output _cvpt_1548;   // oc8051_tb.v(104)
    output _cvpt_1549;   // oc8051_tb.v(104)
    output _cvpt_1550;   // oc8051_tb.v(104)
    output _cvpt_1551;   // oc8051_tb.v(104)
    output _cvpt_1552;   // oc8051_tb.v(104)
    output _cvpt_1553;   // oc8051_tb.v(104)
    output _cvpt_1554;   // oc8051_tb.v(104)
    output _cvpt_1555;   // oc8051_tb.v(104)
    output _cvpt_1556;   // oc8051_tb.v(104)
    output _cvpt_1557;   // oc8051_tb.v(104)
    output _cvpt_1558;   // oc8051_tb.v(104)
    output _cvpt_1559;   // oc8051_tb.v(104)
    output _cvpt_1560;   // oc8051_tb.v(104)
    output _cvpt_1561;   // oc8051_tb.v(104)
    output _cvpt_1562;   // oc8051_tb.v(104)
    output _cvpt_1563;   // oc8051_tb.v(104)
    output _cvpt_1564;   // oc8051_tb.v(104)
    output _cvpt_1565;   // oc8051_tb.v(104)
    output _cvpt_1566;   // oc8051_tb.v(104)
    output _cvpt_1567;   // oc8051_tb.v(104)
    output _cvpt_1568;   // oc8051_tb.v(104)
    output _cvpt_1569;   // oc8051_tb.v(104)
    output _cvpt_1570;   // oc8051_tb.v(104)
    output _cvpt_1571;   // oc8051_tb.v(104)
    output _cvpt_1572;   // oc8051_tb.v(104)
    output _cvpt_1573;   // oc8051_tb.v(104)
    output _cvpt_1574;   // oc8051_tb.v(104)
    output _cvpt_1575;   // oc8051_tb.v(104)
    output _cvpt_1576;   // oc8051_tb.v(104)
    output _cvpt_1577;   // oc8051_tb.v(104)
    output _cvpt_1578;   // oc8051_tb.v(104)
    output _cvpt_1579;   // oc8051_tb.v(104)
    output _cvpt_1580;   // oc8051_tb.v(104)
    output _cvpt_1581;   // oc8051_tb.v(104)
    output _cvpt_1582;   // oc8051_tb.v(104)
    output _cvpt_1583;   // oc8051_tb.v(104)
    output _cvpt_1584;   // oc8051_tb.v(104)
    output _cvpt_1585;   // oc8051_tb.v(104)
    output _cvpt_1586;   // oc8051_tb.v(104)
    output _cvpt_1587;   // oc8051_tb.v(104)
    output _cvpt_1588;   // oc8051_tb.v(104)
    output _cvpt_1589;   // oc8051_tb.v(104)
    output _cvpt_1590;   // oc8051_tb.v(104)
    output _cvpt_1591;   // oc8051_tb.v(104)
    output _cvpt_1592;   // oc8051_tb.v(104)
    output _cvpt_1593;   // oc8051_tb.v(104)
    output _cvpt_1594;   // oc8051_tb.v(104)
    output _cvpt_1595;   // oc8051_tb.v(104)
    output _cvpt_1596;   // oc8051_tb.v(104)
    output _cvpt_1597;   // oc8051_tb.v(104)
    output _cvpt_1598;   // oc8051_tb.v(104)
    output _cvpt_1599;   // oc8051_tb.v(104)
    output _cvpt_1600;   // oc8051_tb.v(104)
    output _cvpt_1601;   // oc8051_tb.v(104)
    output _cvpt_1602;   // oc8051_tb.v(104)
    output _cvpt_1603;   // oc8051_tb.v(104)
    output _cvpt_1604;   // oc8051_tb.v(104)
    output _cvpt_1605;   // oc8051_tb.v(104)
    output _cvpt_1606;   // oc8051_tb.v(104)
    output _cvpt_1607;   // oc8051_tb.v(104)
    output _cvpt_1608;   // oc8051_tb.v(104)
    output _cvpt_1609;   // oc8051_tb.v(104)
    output _cvpt_1610;   // oc8051_tb.v(104)
    output _cvpt_1611;   // oc8051_tb.v(104)
    output _cvpt_1612;   // oc8051_tb.v(104)
    output _cvpt_1613;   // oc8051_tb.v(104)
    output _cvpt_1614;   // oc8051_tb.v(104)
    output _cvpt_1615;   // oc8051_tb.v(104)
    output _cvpt_1616;   // oc8051_tb.v(104)
    output _cvpt_1617;   // oc8051_tb.v(104)
    output _cvpt_1618;   // oc8051_tb.v(104)
    output _cvpt_1619;   // oc8051_tb.v(104)
    output _cvpt_1620;   // oc8051_tb.v(104)
    output _cvpt_1621;   // oc8051_tb.v(104)
    output _cvpt_1622;   // oc8051_tb.v(104)
    output _cvpt_1623;   // oc8051_tb.v(104)
    output _cvpt_1624;   // oc8051_tb.v(104)
    output _cvpt_1625;   // oc8051_tb.v(104)
    output _cvpt_1626;   // oc8051_tb.v(104)
    output _cvpt_1627;   // oc8051_tb.v(104)
    output _cvpt_1628;   // oc8051_tb.v(104)
    output _cvpt_1629;   // oc8051_tb.v(104)
    output _cvpt_1630;   // oc8051_tb.v(104)
    output _cvpt_1631;   // oc8051_tb.v(104)
    output _cvpt_1632;   // oc8051_tb.v(104)
    output _cvpt_1633;   // oc8051_tb.v(104)
    output _cvpt_1634;   // oc8051_tb.v(104)
    output _cvpt_1635;   // oc8051_tb.v(104)
    output _cvpt_1636;   // oc8051_tb.v(104)
    output _cvpt_1637;   // oc8051_tb.v(104)
    output _cvpt_1638;   // oc8051_tb.v(104)
    output _cvpt_1639;   // oc8051_tb.v(104)
    output _cvpt_1640;   // oc8051_tb.v(104)
    output _cvpt_1641;   // oc8051_tb.v(104)
    output _cvpt_1642;   // oc8051_tb.v(104)
    output _cvpt_1643;   // oc8051_tb.v(104)
    output _cvpt_1644;   // oc8051_tb.v(104)
    output _cvpt_1645;   // oc8051_tb.v(104)
    output _cvpt_1646;   // oc8051_tb.v(104)
    output _cvpt_1647;   // oc8051_tb.v(104)
    output _cvpt_1648;   // oc8051_tb.v(104)
    output _cvpt_1649;   // oc8051_tb.v(104)
    output _cvpt_1650;   // oc8051_tb.v(104)
    output _cvpt_1651;   // oc8051_tb.v(104)
    output _cvpt_1652;   // oc8051_tb.v(104)
    output _cvpt_1653;   // oc8051_tb.v(104)
    output _cvpt_1654;   // oc8051_tb.v(104)
    output _cvpt_1655;   // oc8051_tb.v(104)
    output _cvpt_1656;   // oc8051_tb.v(104)
    output _cvpt_1657;   // oc8051_tb.v(104)
    output _cvpt_1658;   // oc8051_tb.v(104)
    output _cvpt_1659;   // oc8051_tb.v(104)
    output _cvpt_1660;   // oc8051_tb.v(104)
    output _cvpt_1661;   // oc8051_tb.v(104)
    output _cvpt_1662;   // oc8051_tb.v(104)
    output _cvpt_1663;   // oc8051_tb.v(104)
    output _cvpt_1664;   // oc8051_tb.v(104)
    output _cvpt_1665;   // oc8051_tb.v(104)
    output _cvpt_1666;   // oc8051_tb.v(104)
    output _cvpt_1667;   // oc8051_tb.v(104)
    output _cvpt_1668;   // oc8051_tb.v(104)
    output _cvpt_1669;   // oc8051_tb.v(104)
    output _cvpt_1670;   // oc8051_tb.v(104)
    output _cvpt_1671;   // oc8051_tb.v(104)
    output _cvpt_1672;   // oc8051_tb.v(104)
    output _cvpt_1673;   // oc8051_tb.v(104)
    output _cvpt_1674;   // oc8051_tb.v(104)
    output _cvpt_1675;   // oc8051_tb.v(104)
    output _cvpt_1676;   // oc8051_tb.v(104)
    output _cvpt_1677;   // oc8051_tb.v(104)
    output _cvpt_1678;   // oc8051_tb.v(104)
    output _cvpt_1679;   // oc8051_tb.v(104)
    output _cvpt_1680;   // oc8051_tb.v(104)
    output _cvpt_1681;   // oc8051_tb.v(104)
    output _cvpt_1682;   // oc8051_tb.v(104)
    output _cvpt_1683;   // oc8051_tb.v(104)
    output _cvpt_1684;   // oc8051_tb.v(104)
    output _cvpt_1685;   // oc8051_tb.v(104)
    output _cvpt_1686;   // oc8051_tb.v(104)
    output _cvpt_1687;   // oc8051_tb.v(104)
    output _cvpt_1688;   // oc8051_tb.v(104)
    output _cvpt_1689;   // oc8051_tb.v(104)
    output _cvpt_1690;   // oc8051_tb.v(104)
    output _cvpt_1691;   // oc8051_tb.v(104)
    output _cvpt_1692;   // oc8051_tb.v(104)
    output _cvpt_1693;   // oc8051_tb.v(104)
    output _cvpt_1694;   // oc8051_tb.v(104)
    output _cvpt_1695;   // oc8051_tb.v(104)
    output _cvpt_1696;   // oc8051_tb.v(104)
    output _cvpt_1697;   // oc8051_tb.v(104)
    output _cvpt_1698;   // oc8051_tb.v(104)
    output _cvpt_1699;   // oc8051_tb.v(104)
    output _cvpt_1700;   // oc8051_tb.v(104)
    output _cvpt_1701;   // oc8051_tb.v(104)
    output _cvpt_1702;   // oc8051_tb.v(104)
    output _cvpt_1703;   // oc8051_tb.v(104)
    output _cvpt_1704;   // oc8051_tb.v(104)
    output _cvpt_1705;   // oc8051_tb.v(104)
    output _cvpt_1706;   // oc8051_tb.v(104)
    output _cvpt_1707;   // oc8051_tb.v(104)
    output _cvpt_1708;   // oc8051_tb.v(104)
    output _cvpt_1709;   // oc8051_tb.v(104)
    output _cvpt_1710;   // oc8051_tb.v(104)
    output _cvpt_1711;   // oc8051_tb.v(104)
    output _cvpt_1712;   // oc8051_tb.v(104)
    output _cvpt_1713;   // oc8051_tb.v(104)
    output _cvpt_1714;   // oc8051_tb.v(104)
    output _cvpt_1715;   // oc8051_tb.v(104)
    output _cvpt_1716;   // oc8051_tb.v(104)
    output _cvpt_1717;   // oc8051_tb.v(104)
    output _cvpt_1718;   // oc8051_tb.v(104)
    output _cvpt_1719;   // oc8051_tb.v(104)
    output _cvpt_1720;   // oc8051_tb.v(104)
    output _cvpt_1721;   // oc8051_tb.v(104)
    output _cvpt_1722;   // oc8051_tb.v(104)
    output _cvpt_1723;   // oc8051_tb.v(104)
    output _cvpt_1724;   // oc8051_tb.v(104)
    output _cvpt_1725;   // oc8051_tb.v(104)
    output _cvpt_1726;   // oc8051_tb.v(104)
    output _cvpt_1727;   // oc8051_tb.v(104)
    output _cvpt_1728;   // oc8051_tb.v(104)
    output _cvpt_1729;   // oc8051_tb.v(104)
    output _cvpt_1730;   // oc8051_tb.v(104)
    output _cvpt_1731;   // oc8051_tb.v(104)
    output _cvpt_1732;   // oc8051_tb.v(104)
    output _cvpt_1733;   // oc8051_tb.v(104)
    output _cvpt_1734;   // oc8051_tb.v(104)
    output _cvpt_1735;   // oc8051_tb.v(104)
    output _cvpt_1736;   // oc8051_tb.v(104)
    output _cvpt_1737;   // oc8051_tb.v(104)
    output _cvpt_1738;   // oc8051_tb.v(104)
    output _cvpt_1739;   // oc8051_tb.v(104)
    output _cvpt_1740;   // oc8051_tb.v(104)
    output _cvpt_1741;   // oc8051_tb.v(104)
    output _cvpt_1742;   // oc8051_tb.v(104)
    output _cvpt_1743;   // oc8051_tb.v(104)
    output _cvpt_1744;   // oc8051_tb.v(104)
    output _cvpt_1745;   // oc8051_tb.v(104)
    output _cvpt_1746;   // oc8051_tb.v(104)
    output _cvpt_1747;   // oc8051_tb.v(104)
    output _cvpt_1748;   // oc8051_tb.v(104)
    output _cvpt_1749;   // oc8051_tb.v(104)
    output _cvpt_1750;   // oc8051_tb.v(104)
    output _cvpt_1751;   // oc8051_tb.v(104)
    output _cvpt_1752;   // oc8051_tb.v(104)
    output _cvpt_1753;   // oc8051_tb.v(104)
    output _cvpt_1754;   // oc8051_tb.v(104)
    output _cvpt_1755;   // oc8051_tb.v(104)
    output _cvpt_1756;   // oc8051_tb.v(104)
    output _cvpt_1757;   // oc8051_tb.v(104)
    output _cvpt_1758;   // oc8051_tb.v(104)
    output _cvpt_1759;   // oc8051_tb.v(104)
    output _cvpt_1760;   // oc8051_tb.v(104)
    output _cvpt_1761;   // oc8051_tb.v(104)
    output _cvpt_1762;   // oc8051_tb.v(104)
    output _cvpt_1763;   // oc8051_tb.v(104)
    output _cvpt_1764;   // oc8051_tb.v(104)
    output _cvpt_1765;   // oc8051_tb.v(104)
    output _cvpt_1766;   // oc8051_tb.v(104)
    output _cvpt_1767;   // oc8051_tb.v(104)
    output _cvpt_1768;   // oc8051_tb.v(104)
    output _cvpt_1769;   // oc8051_tb.v(104)
    output _cvpt_1770;   // oc8051_tb.v(104)
    output _cvpt_1771;   // oc8051_tb.v(104)
    output _cvpt_1772;   // oc8051_tb.v(104)
    output _cvpt_1773;   // oc8051_tb.v(104)
    output _cvpt_1774;   // oc8051_tb.v(104)
    output _cvpt_1775;   // oc8051_tb.v(104)
    output _cvpt_1776;   // oc8051_tb.v(104)
    output _cvpt_1777;   // oc8051_tb.v(104)
    output _cvpt_1778;   // oc8051_tb.v(104)
    output _cvpt_1779;   // oc8051_tb.v(104)
    output _cvpt_1780;   // oc8051_tb.v(104)
    output _cvpt_1781;   // oc8051_tb.v(104)
    output _cvpt_1782;   // oc8051_tb.v(104)
    output _cvpt_1783;   // oc8051_tb.v(104)
    output _cvpt_1784;   // oc8051_tb.v(104)
    output _cvpt_1785;   // oc8051_tb.v(104)
    output _cvpt_1786;   // oc8051_tb.v(104)
    output _cvpt_1787;   // oc8051_tb.v(104)
    output _cvpt_1788;   // oc8051_tb.v(104)
    output _cvpt_1789;   // oc8051_tb.v(104)
    output _cvpt_1790;   // oc8051_tb.v(104)
    output _cvpt_1791;   // oc8051_tb.v(104)
    output _cvpt_1792;   // oc8051_tb.v(104)
    output _cvpt_1793;   // oc8051_tb.v(104)
    output _cvpt_1794;   // oc8051_tb.v(104)
    output _cvpt_1795;   // oc8051_tb.v(104)
    output _cvpt_1796;   // oc8051_tb.v(104)
    output _cvpt_1797;   // oc8051_tb.v(104)
    output _cvpt_1798;   // oc8051_tb.v(104)
    output _cvpt_1799;   // oc8051_tb.v(104)
    output _cvpt_1800;   // oc8051_tb.v(104)
    output _cvpt_1801;   // oc8051_tb.v(104)
    output _cvpt_1802;   // oc8051_tb.v(104)
    output _cvpt_1803;   // oc8051_tb.v(104)
    output _cvpt_1804;   // oc8051_tb.v(104)
    output _cvpt_1805;   // oc8051_tb.v(104)
    output _cvpt_1806;   // oc8051_tb.v(104)
    output _cvpt_1807;   // oc8051_tb.v(104)
    output _cvpt_1808;   // oc8051_tb.v(104)
    output _cvpt_1809;   // oc8051_tb.v(104)
    output _cvpt_1810;   // oc8051_tb.v(104)
    output _cvpt_1811;   // oc8051_tb.v(104)
    output _cvpt_1812;   // oc8051_tb.v(104)
    output _cvpt_1813;   // oc8051_tb.v(104)
    output _cvpt_1814;   // oc8051_tb.v(104)
    output _cvpt_1815;   // oc8051_tb.v(104)
    output _cvpt_1816;   // oc8051_tb.v(104)
    output _cvpt_1817;   // oc8051_tb.v(104)
    output _cvpt_1818;   // oc8051_tb.v(104)
    output _cvpt_1819;   // oc8051_tb.v(104)
    output _cvpt_1820;   // oc8051_tb.v(104)
    output _cvpt_1821;   // oc8051_tb.v(104)
    output _cvpt_1822;   // oc8051_tb.v(104)
    output _cvpt_1823;   // oc8051_tb.v(104)
    output _cvpt_1824;   // oc8051_tb.v(104)
    output _cvpt_1825;   // oc8051_tb.v(104)
    output _cvpt_1826;   // oc8051_tb.v(104)
    output _cvpt_1827;   // oc8051_tb.v(104)
    output _cvpt_1828;   // oc8051_tb.v(104)
    output _cvpt_1829;   // oc8051_tb.v(104)
    output _cvpt_1830;   // oc8051_tb.v(104)
    output _cvpt_1831;   // oc8051_tb.v(104)
    output _cvpt_1832;   // oc8051_tb.v(104)
    output _cvpt_1833;   // oc8051_tb.v(104)
    output _cvpt_1834;   // oc8051_tb.v(104)
    output _cvpt_1835;   // oc8051_tb.v(104)
    output _cvpt_1836;   // oc8051_tb.v(104)
    output _cvpt_1837;   // oc8051_tb.v(104)
    output _cvpt_1838;   // oc8051_tb.v(104)
    output _cvpt_1839;   // oc8051_tb.v(104)
    output _cvpt_1840;   // oc8051_tb.v(104)
    output _cvpt_1841;   // oc8051_tb.v(104)
    output _cvpt_1842;   // oc8051_tb.v(104)
    output _cvpt_1843;   // oc8051_tb.v(104)
    output _cvpt_1844;   // oc8051_tb.v(104)
    output _cvpt_1845;   // oc8051_tb.v(104)
    output _cvpt_1846;   // oc8051_tb.v(104)
    output _cvpt_1847;   // oc8051_tb.v(104)
    output _cvpt_1848;   // oc8051_tb.v(104)
    output _cvpt_1849;   // oc8051_tb.v(104)
    output _cvpt_1850;   // oc8051_tb.v(104)
    output _cvpt_1851;   // oc8051_tb.v(104)
    output _cvpt_1852;   // oc8051_tb.v(104)
    output _cvpt_1853;   // oc8051_tb.v(104)
    output _cvpt_1854;   // oc8051_tb.v(104)
    output _cvpt_1855;   // oc8051_tb.v(104)
    output _cvpt_1856;   // oc8051_tb.v(104)
    output _cvpt_1857;   // oc8051_tb.v(104)
    output _cvpt_1858;   // oc8051_tb.v(104)
    output _cvpt_1859;   // oc8051_tb.v(104)
    output _cvpt_1860;   // oc8051_tb.v(104)
    output _cvpt_1861;   // oc8051_tb.v(104)
    output _cvpt_1862;   // oc8051_tb.v(104)
    output _cvpt_1863;   // oc8051_tb.v(104)
    output _cvpt_1864;   // oc8051_tb.v(104)
    output _cvpt_1865;   // oc8051_tb.v(104)
    output _cvpt_1866;   // oc8051_tb.v(104)
    output _cvpt_1867;   // oc8051_tb.v(104)
    output _cvpt_1868;   // oc8051_tb.v(104)
    output _cvpt_1869;   // oc8051_tb.v(104)
    output _cvpt_1870;   // oc8051_tb.v(104)
    output _cvpt_1871;   // oc8051_tb.v(104)
    output _cvpt_1872;   // oc8051_tb.v(104)
    output _cvpt_1873;   // oc8051_tb.v(104)
    output _cvpt_1874;   // oc8051_tb.v(104)
    output _cvpt_1875;   // oc8051_tb.v(104)
    output _cvpt_1876;   // oc8051_tb.v(104)
    output _cvpt_1877;   // oc8051_tb.v(104)
    output _cvpt_1878;   // oc8051_tb.v(104)
    output _cvpt_1879;   // oc8051_tb.v(104)
    output _cvpt_1880;   // oc8051_tb.v(104)
    output _cvpt_1881;   // oc8051_tb.v(104)
    output _cvpt_1882;   // oc8051_tb.v(104)
    output _cvpt_1883;   // oc8051_tb.v(104)
    output _cvpt_1884;   // oc8051_tb.v(104)
    output _cvpt_1885;   // oc8051_tb.v(104)
    output _cvpt_1886;   // oc8051_tb.v(104)
    output _cvpt_1887;   // oc8051_tb.v(104)
    output _cvpt_1888;   // oc8051_tb.v(104)
    output _cvpt_1889;   // oc8051_tb.v(104)
    output _cvpt_1890;   // oc8051_tb.v(104)
    output _cvpt_1891;   // oc8051_tb.v(104)
    output _cvpt_1892;   // oc8051_tb.v(104)
    output _cvpt_1893;   // oc8051_tb.v(104)
    output _cvpt_1894;   // oc8051_tb.v(104)
    output _cvpt_1895;   // oc8051_tb.v(104)
    output _cvpt_1896;   // oc8051_tb.v(104)
    output _cvpt_1897;   // oc8051_tb.v(104)
    output _cvpt_1898;   // oc8051_tb.v(104)
    output _cvpt_1899;   // oc8051_tb.v(104)
    output _cvpt_1900;   // oc8051_tb.v(104)
    output _cvpt_1901;   // oc8051_tb.v(104)
    output _cvpt_1902;   // oc8051_tb.v(104)
    output _cvpt_1903;   // oc8051_tb.v(104)
    output _cvpt_1904;   // oc8051_tb.v(104)
    output _cvpt_1905;   // oc8051_tb.v(104)
    output _cvpt_1906;   // oc8051_tb.v(104)
    output _cvpt_1907;   // oc8051_tb.v(104)
    output _cvpt_1908;   // oc8051_tb.v(104)
    output _cvpt_1909;   // oc8051_tb.v(104)
    output _cvpt_1910;   // oc8051_tb.v(104)
    output _cvpt_1911;   // oc8051_tb.v(104)
    output _cvpt_1912;   // oc8051_tb.v(104)
    output _cvpt_1913;   // oc8051_tb.v(104)
    output _cvpt_1914;   // oc8051_tb.v(104)
    output _cvpt_1915;   // oc8051_tb.v(104)
    output _cvpt_1916;   // oc8051_tb.v(104)
    output _cvpt_1917;   // oc8051_tb.v(104)
    output _cvpt_1918;   // oc8051_tb.v(104)
    output _cvpt_1919;   // oc8051_tb.v(104)
    output _cvpt_1920;   // oc8051_tb.v(104)
    output _cvpt_1921;   // oc8051_tb.v(104)
    output _cvpt_1922;   // oc8051_tb.v(104)
    output _cvpt_1923;   // oc8051_tb.v(104)
    output _cvpt_1924;   // oc8051_tb.v(104)
    output _cvpt_1925;   // oc8051_tb.v(104)
    output _cvpt_1926;   // oc8051_tb.v(104)
    output _cvpt_1927;   // oc8051_tb.v(104)
    output _cvpt_1928;   // oc8051_tb.v(104)
    output _cvpt_1929;   // oc8051_tb.v(104)
    output _cvpt_1930;   // oc8051_tb.v(104)
    output _cvpt_1931;   // oc8051_tb.v(104)
    output _cvpt_1932;   // oc8051_tb.v(104)
    output _cvpt_1933;   // oc8051_tb.v(104)
    output _cvpt_1934;   // oc8051_tb.v(104)
    output _cvpt_1935;   // oc8051_tb.v(104)
    output _cvpt_1936;   // oc8051_tb.v(104)
    output _cvpt_1937;   // oc8051_tb.v(104)
    output _cvpt_1938;   // oc8051_tb.v(104)
    output _cvpt_1939;   // oc8051_tb.v(104)
    output _cvpt_1940;   // oc8051_tb.v(104)
    output _cvpt_1941;   // oc8051_tb.v(104)
    output _cvpt_1942;   // oc8051_tb.v(104)
    output _cvpt_1943;   // oc8051_tb.v(104)
    output _cvpt_1944;   // oc8051_tb.v(104)
    output _cvpt_1945;   // oc8051_tb.v(104)
    output _cvpt_1946;   // oc8051_tb.v(104)
    output _cvpt_1947;   // oc8051_tb.v(104)
    output _cvpt_1948;   // oc8051_tb.v(104)
    output _cvpt_1949;   // oc8051_tb.v(104)
    output _cvpt_1950;   // oc8051_tb.v(104)
    output _cvpt_1951;   // oc8051_tb.v(104)
    output _cvpt_1952;   // oc8051_tb.v(104)
    output _cvpt_1953;   // oc8051_tb.v(104)
    output _cvpt_1954;   // oc8051_tb.v(104)
    output _cvpt_1955;   // oc8051_tb.v(104)
    output _cvpt_1956;   // oc8051_tb.v(104)
    output _cvpt_1957;   // oc8051_tb.v(104)
    output _cvpt_1958;   // oc8051_tb.v(104)
    output _cvpt_1959;   // oc8051_tb.v(104)
    output _cvpt_1960;   // oc8051_tb.v(104)
    output _cvpt_1961;   // oc8051_tb.v(104)
    output _cvpt_1962;   // oc8051_tb.v(104)
    output _cvpt_1963;   // oc8051_tb.v(104)
    output _cvpt_1964;   // oc8051_tb.v(104)
    output _cvpt_1965;   // oc8051_tb.v(104)
    output _cvpt_1966;   // oc8051_tb.v(104)
    output _cvpt_1967;   // oc8051_tb.v(104)
    output _cvpt_1968;   // oc8051_tb.v(104)
    output _cvpt_1969;   // oc8051_tb.v(104)
    output _cvpt_1970;   // oc8051_tb.v(104)
    output _cvpt_1971;   // oc8051_tb.v(104)
    output _cvpt_1972;   // oc8051_tb.v(104)
    output _cvpt_1973;   // oc8051_tb.v(104)
    output _cvpt_1974;   // oc8051_tb.v(104)
    output _cvpt_1975;   // oc8051_tb.v(104)
    output _cvpt_1976;   // oc8051_tb.v(104)
    output _cvpt_1977;   // oc8051_tb.v(104)
    output _cvpt_1978;   // oc8051_tb.v(104)
    output _cvpt_1979;   // oc8051_tb.v(104)
    output _cvpt_1980;   // oc8051_tb.v(104)
    output _cvpt_1981;   // oc8051_tb.v(104)
    output _cvpt_1982;   // oc8051_tb.v(104)
    output _cvpt_1983;   // oc8051_tb.v(104)
    output _cvpt_1984;   // oc8051_tb.v(104)
    output _cvpt_1985;   // oc8051_tb.v(104)
    output _cvpt_1986;   // oc8051_tb.v(104)
    output _cvpt_1987;   // oc8051_tb.v(104)
    output _cvpt_1988;   // oc8051_tb.v(104)
    output _cvpt_1989;   // oc8051_tb.v(104)
    output _cvpt_1990;   // oc8051_tb.v(104)
    output _cvpt_1991;   // oc8051_tb.v(104)
    output _cvpt_1992;   // oc8051_tb.v(104)
    output _cvpt_1993;   // oc8051_tb.v(104)
    output _cvpt_1994;   // oc8051_tb.v(104)
    output _cvpt_1995;   // oc8051_tb.v(104)
    output _cvpt_1996;   // oc8051_tb.v(104)
    output _cvpt_1997;   // oc8051_tb.v(104)
    output _cvpt_1998;   // oc8051_tb.v(104)
    output _cvpt_1999;   // oc8051_tb.v(104)
    output _cvpt_2000;   // oc8051_tb.v(104)
    output _cvpt_2001;   // oc8051_tb.v(104)
    output _cvpt_2002;   // oc8051_tb.v(104)
    output _cvpt_2003;   // oc8051_tb.v(104)
    output _cvpt_2004;   // oc8051_tb.v(104)
    output _cvpt_2005;   // oc8051_tb.v(104)
    output _cvpt_2006;   // oc8051_tb.v(104)
    output _cvpt_2007;   // oc8051_tb.v(104)
    output _cvpt_2008;   // oc8051_tb.v(104)
    output _cvpt_2009;   // oc8051_tb.v(104)
    output _cvpt_2010;   // oc8051_tb.v(104)
    output _cvpt_2011;   // oc8051_tb.v(104)
    output _cvpt_2012;   // oc8051_tb.v(104)
    output _cvpt_2013;   // oc8051_tb.v(104)
    output _cvpt_2014;   // oc8051_tb.v(104)
    output _cvpt_2015;   // oc8051_tb.v(104)
    output _cvpt_2016;   // oc8051_tb.v(104)
    output _cvpt_2017;   // oc8051_tb.v(104)
    output _cvpt_2018;   // oc8051_tb.v(104)
    output _cvpt_2019;   // oc8051_tb.v(104)
    output _cvpt_2020;   // oc8051_tb.v(104)
    output _cvpt_2021;   // oc8051_tb.v(104)
    output _cvpt_2022;   // oc8051_tb.v(104)
    output _cvpt_2023;   // oc8051_tb.v(104)
    output _cvpt_2024;   // oc8051_tb.v(104)
    output _cvpt_2025;   // oc8051_tb.v(104)
    output _cvpt_2026;   // oc8051_tb.v(104)
    output _cvpt_2027;   // oc8051_tb.v(104)
    output _cvpt_2028;   // oc8051_tb.v(104)
    output _cvpt_2029;   // oc8051_tb.v(104)
    output _cvpt_2030;   // oc8051_tb.v(104)
    output _cvpt_2031;   // oc8051_tb.v(104)
    output _cvpt_2032;   // oc8051_tb.v(104)
    output _cvpt_2033;   // oc8051_tb.v(104)
    output _cvpt_2034;   // oc8051_tb.v(104)
    output _cvpt_2035;   // oc8051_tb.v(104)
    output _cvpt_2036;   // oc8051_tb.v(104)
    output _cvpt_2037;   // oc8051_tb.v(104)
    output _cvpt_2038;   // oc8051_tb.v(104)
    output _cvpt_2039;   // oc8051_tb.v(104)
    output _cvpt_2040;   // oc8051_tb.v(104)
    output _cvpt_2041;   // oc8051_tb.v(104)
    output _cvpt_2042;   // oc8051_tb.v(104)
    output _cvpt_2043;   // oc8051_tb.v(104)
    output _cvpt_2044;   // oc8051_tb.v(104)
    output _cvpt_2045;   // oc8051_tb.v(104)
    output _cvpt_2046;   // oc8051_tb.v(104)
    output _cvpt_2047;   // oc8051_tb.v(104)
    output _cvpt_2048;   // oc8051_tb.v(104)
    output _cvpt_2049;   // oc8051_tb.v(104)
    output _cvpt_2050;   // oc8051_tb.v(104)
    output _cvpt_2051;   // oc8051_tb.v(104)
    output _cvpt_2052;   // oc8051_tb.v(104)
    output _cvpt_2053;   // oc8051_tb.v(104)
    output _cvpt_2054;   // oc8051_tb.v(104)
    output _cvpt_2055;   // oc8051_tb.v(104)
    output _cvpt_2056;   // oc8051_tb.v(104)
    output _cvpt_2057;   // oc8051_tb.v(104)
    output _cvpt_2058;   // oc8051_tb.v(104)
    output _cvpt_2059;   // oc8051_tb.v(104)
    output _cvpt_2060;   // oc8051_tb.v(104)
    output _cvpt_2061;   // oc8051_tb.v(104)
    output _cvpt_2062;   // oc8051_tb.v(104)
    output _cvpt_2063;   // oc8051_tb.v(104)
    output _cvpt_2064;   // oc8051_tb.v(104)
    output _cvpt_2065;   // oc8051_tb.v(104)
    output _cvpt_2066;   // oc8051_tb.v(104)
    output _cvpt_2067;   // oc8051_tb.v(104)
    output _cvpt_2068;   // oc8051_tb.v(104)
    output _cvpt_2069;   // oc8051_tb.v(104)
    output _cvpt_2070;   // oc8051_tb.v(104)
    output _cvpt_2071;   // oc8051_tb.v(104)
    output _cvpt_2072;   // oc8051_tb.v(104)
    output _cvpt_2073;   // oc8051_tb.v(104)
    output _cvpt_2074;   // oc8051_tb.v(104)
    output _cvpt_2075;   // oc8051_tb.v(104)
    output _cvpt_2076;   // oc8051_tb.v(104)
    output _cvpt_2077;   // oc8051_tb.v(104)
    output _cvpt_2078;   // oc8051_tb.v(104)
    output _cvpt_2079;   // oc8051_tb.v(104)
    output _cvpt_2080;   // oc8051_tb.v(104)
    output _cvpt_2081;   // oc8051_tb.v(104)
    output _cvpt_2082;   // oc8051_tb.v(104)
    output _cvpt_2083;   // oc8051_tb.v(104)
    output _cvpt_2084;   // oc8051_tb.v(104)
    output _cvpt_2085;   // oc8051_tb.v(104)
    output _cvpt_2086;   // oc8051_tb.v(104)
    output _cvpt_2087;   // oc8051_tb.v(104)
    output _cvpt_2088;   // oc8051_tb.v(104)
    output _cvpt_2089;   // oc8051_tb.v(104)
    output _cvpt_2090;   // oc8051_tb.v(104)
    output _cvpt_2091;   // oc8051_tb.v(104)
    output _cvpt_2092;   // oc8051_tb.v(104)
    output _cvpt_2093;   // oc8051_tb.v(104)
    output _cvpt_2094;   // oc8051_tb.v(104)
    output _cvpt_2095;   // oc8051_tb.v(104)
    output _cvpt_2096;   // oc8051_tb.v(104)
    output _cvpt_2097;   // oc8051_tb.v(104)
    output _cvpt_2098;   // oc8051_tb.v(104)
    output _cvpt_2099;   // oc8051_tb.v(104)
    output _cvpt_2100;   // oc8051_tb.v(104)
    output _cvpt_2101;   // oc8051_tb.v(104)
    output _cvpt_2102;   // oc8051_tb.v(104)
    output _cvpt_2103;   // oc8051_tb.v(104)
    output _cvpt_2104;   // oc8051_tb.v(104)
    output _cvpt_2105;   // oc8051_tb.v(104)
    output _cvpt_2106;   // oc8051_tb.v(104)
    output _cvpt_2107;   // oc8051_tb.v(104)
    output _cvpt_2108;   // oc8051_tb.v(104)
    output _cvpt_2109;   // oc8051_tb.v(104)
    output _cvpt_2110;   // oc8051_tb.v(104)
    output _cvpt_2111;   // oc8051_tb.v(104)
    output _cvpt_2112;   // oc8051_tb.v(104)
    output _cvpt_2113;   // oc8051_tb.v(104)
    output _cvpt_2114;   // oc8051_tb.v(104)
    output _cvpt_2115;   // oc8051_tb.v(104)
    output _cvpt_2116;   // oc8051_tb.v(104)
    output _cvpt_2117;   // oc8051_tb.v(104)
    output _cvpt_2118;   // oc8051_tb.v(104)
    output _cvpt_2119;   // oc8051_tb.v(104)
    output _cvpt_2120;   // oc8051_tb.v(104)
    output _cvpt_2121;   // oc8051_tb.v(104)
    output _cvpt_2122;   // oc8051_tb.v(104)
    output _cvpt_2123;   // oc8051_tb.v(104)
    output _cvpt_2124;   // oc8051_tb.v(104)
    output _cvpt_2125;   // oc8051_tb.v(104)
    output _cvpt_2126;   // oc8051_tb.v(104)
    output _cvpt_2127;   // oc8051_tb.v(104)
    output _cvpt_2128;   // oc8051_tb.v(104)
    output _cvpt_2129;   // oc8051_tb.v(104)
    output _cvpt_2130;   // oc8051_tb.v(104)
    output _cvpt_2131;   // oc8051_tb.v(104)
    output _cvpt_2132;   // oc8051_tb.v(104)
    output _cvpt_2133;   // oc8051_tb.v(104)
    output _cvpt_2134;   // oc8051_tb.v(104)
    output _cvpt_2135;   // oc8051_tb.v(104)
    output _cvpt_2136;   // oc8051_tb.v(104)
    output _cvpt_2137;   // oc8051_tb.v(104)
    output _cvpt_2138;   // oc8051_tb.v(104)
    output _cvpt_2139;   // oc8051_tb.v(104)
    output _cvpt_2140;   // oc8051_tb.v(104)
    output _cvpt_2141;   // oc8051_tb.v(104)
    output _cvpt_2142;   // oc8051_tb.v(104)
    output _cvpt_2143;   // oc8051_tb.v(104)
    output _cvpt_2144;   // oc8051_tb.v(104)
    output _cvpt_2145;   // oc8051_tb.v(104)
    output _cvpt_2146;   // oc8051_tb.v(104)
    output _cvpt_2147;   // oc8051_tb.v(104)
    output _cvpt_2148;   // oc8051_tb.v(104)
    output _cvpt_2149;   // oc8051_tb.v(104)
    output _cvpt_2150;   // oc8051_tb.v(104)
    output _cvpt_2151;   // oc8051_tb.v(104)
    output _cvpt_2152;   // oc8051_tb.v(104)
    output _cvpt_2153;   // oc8051_tb.v(104)
    output _cvpt_2154;   // oc8051_tb.v(104)
    output _cvpt_2155;   // oc8051_tb.v(104)
    output _cvpt_2156;   // oc8051_tb.v(104)
    output _cvpt_2157;   // oc8051_tb.v(104)
    output _cvpt_2158;   // oc8051_tb.v(104)
    output _cvpt_2159;   // oc8051_tb.v(104)
    output _cvpt_2160;   // oc8051_tb.v(104)
    output _cvpt_2161;   // oc8051_tb.v(104)
    output _cvpt_2162;   // oc8051_tb.v(104)
    output _cvpt_2163;   // oc8051_tb.v(104)
    output _cvpt_2164;   // oc8051_tb.v(104)
    output _cvpt_2165;   // oc8051_tb.v(104)
    output _cvpt_2166;   // oc8051_tb.v(104)
    output _cvpt_2167;   // oc8051_tb.v(104)
    output _cvpt_2168;   // oc8051_tb.v(104)
    output _cvpt_2169;   // oc8051_tb.v(104)
    output _cvpt_2170;   // oc8051_tb.v(104)
    output _cvpt_2171;   // oc8051_tb.v(104)
    output _cvpt_2172;   // oc8051_tb.v(104)
    output _cvpt_2173;   // oc8051_tb.v(104)
    output _cvpt_2174;   // oc8051_tb.v(104)
    output _cvpt_2175;   // oc8051_tb.v(104)
    output _cvpt_2176;   // oc8051_tb.v(104)
    output _cvpt_2177;   // oc8051_tb.v(104)
    output _cvpt_2178;   // oc8051_tb.v(104)
    output _cvpt_2179;   // oc8051_tb.v(104)
    output _cvpt_2180;   // oc8051_tb.v(104)
    output _cvpt_2181;   // oc8051_tb.v(104)
    output _cvpt_2182;   // oc8051_tb.v(104)
    output _cvpt_2183;   // oc8051_tb.v(104)
    output _cvpt_2184;   // oc8051_tb.v(104)
    output _cvpt_2185;   // oc8051_tb.v(104)
    output _cvpt_2186;   // oc8051_tb.v(104)
    output _cvpt_2187;   // oc8051_tb.v(104)
    output _cvpt_2188;   // oc8051_tb.v(104)
    output _cvpt_2189;   // oc8051_tb.v(104)
    output _cvpt_2190;   // oc8051_tb.v(104)
    output _cvpt_2191;   // oc8051_tb.v(104)
    output _cvpt_2192;   // oc8051_tb.v(104)
    output _cvpt_2193;   // oc8051_tb.v(104)
    output _cvpt_2194;   // oc8051_tb.v(104)
    output _cvpt_2195;   // oc8051_tb.v(104)
    output _cvpt_2196;   // oc8051_tb.v(104)
    output _cvpt_2197;   // oc8051_tb.v(104)
    output _cvpt_2198;   // oc8051_tb.v(104)
    output _cvpt_2199;   // oc8051_tb.v(104)
    output _cvpt_2200;   // oc8051_tb.v(104)
    output _cvpt_2201;   // oc8051_tb.v(104)
    output _cvpt_2202;   // oc8051_tb.v(104)
    output _cvpt_2203;   // oc8051_tb.v(104)
    output _cvpt_2204;   // oc8051_tb.v(104)
    output _cvpt_2205;   // oc8051_tb.v(104)
    output _cvpt_2206;   // oc8051_tb.v(104)
    output _cvpt_2207;   // oc8051_tb.v(104)
    output _cvpt_2208;   // oc8051_tb.v(104)
    output _cvpt_2209;   // oc8051_tb.v(104)
    output _cvpt_2210;   // oc8051_tb.v(104)
    output _cvpt_2211;   // oc8051_tb.v(104)
    output _cvpt_2212;   // oc8051_tb.v(104)
    output _cvpt_2213;   // oc8051_tb.v(104)
    output _cvpt_2214;   // oc8051_tb.v(104)
    output _cvpt_2215;   // oc8051_tb.v(104)
    output _cvpt_2216;   // oc8051_tb.v(104)
    output _cvpt_2217;   // oc8051_tb.v(104)
    output _cvpt_2218;   // oc8051_tb.v(104)
    output _cvpt_2219;   // oc8051_tb.v(104)
    output _cvpt_2220;   // oc8051_tb.v(104)
    output _cvpt_2221;   // oc8051_tb.v(104)
    output _cvpt_2222;   // oc8051_tb.v(104)
    output _cvpt_2223;   // oc8051_tb.v(104)
    output _cvpt_2224;   // oc8051_tb.v(104)
    output _cvpt_2225;   // oc8051_tb.v(104)
    output _cvpt_2226;   // oc8051_tb.v(104)
    output _cvpt_2227;   // oc8051_tb.v(104)
    output _cvpt_2228;   // oc8051_tb.v(104)
    output _cvpt_2229;   // oc8051_tb.v(104)
    output _cvpt_2230;   // oc8051_tb.v(104)
    output _cvpt_2231;   // oc8051_tb.v(104)
    output _cvpt_2232;   // oc8051_tb.v(104)
    output _cvpt_2233;   // oc8051_tb.v(104)
    output _cvpt_2234;   // oc8051_tb.v(104)
    output _cvpt_2235;   // oc8051_tb.v(104)
    output _cvpt_2236;   // oc8051_tb.v(104)
    output _cvpt_2237;   // oc8051_tb.v(104)
    output _cvpt_2238;   // oc8051_tb.v(104)
    output _cvpt_2239;   // oc8051_tb.v(104)
    output _cvpt_2240;   // oc8051_tb.v(104)
    output _cvpt_2241;   // oc8051_tb.v(104)
    output _cvpt_2242;   // oc8051_tb.v(104)
    output _cvpt_2243;   // oc8051_tb.v(104)
    output _cvpt_2244;   // oc8051_tb.v(104)
    output _cvpt_2245;   // oc8051_tb.v(104)
    output _cvpt_2246;   // oc8051_tb.v(104)
    output _cvpt_2247;   // oc8051_tb.v(104)
    output _cvpt_2248;   // oc8051_tb.v(104)
    output _cvpt_2249;   // oc8051_tb.v(104)
    output _cvpt_2250;   // oc8051_tb.v(104)
    output _cvpt_2251;   // oc8051_tb.v(104)
    output _cvpt_2252;   // oc8051_tb.v(104)
    output _cvpt_2253;   // oc8051_tb.v(104)
    output _cvpt_2254;   // oc8051_tb.v(104)
    output _cvpt_2255;   // oc8051_tb.v(104)
    output _cvpt_2256;   // oc8051_tb.v(104)
    output _cvpt_2257;   // oc8051_tb.v(104)
    output _cvpt_2258;   // oc8051_tb.v(104)
    output _cvpt_2259;   // oc8051_tb.v(104)
    output _cvpt_2260;   // oc8051_tb.v(104)
    output _cvpt_2261;   // oc8051_tb.v(104)
    output _cvpt_2262;   // oc8051_tb.v(104)
    output _cvpt_2263;   // oc8051_tb.v(104)
    output _cvpt_2264;   // oc8051_tb.v(104)
    output _cvpt_2265;   // oc8051_tb.v(104)
    output _cvpt_2266;   // oc8051_tb.v(104)
    output _cvpt_2267;   // oc8051_tb.v(104)
    output _cvpt_2268;   // oc8051_tb.v(104)
    output _cvpt_2269;   // oc8051_tb.v(104)
    output _cvpt_2270;   // oc8051_tb.v(104)
    output _cvpt_2271;   // oc8051_tb.v(104)
    output _cvpt_2272;   // oc8051_tb.v(104)
    output _cvpt_2273;   // oc8051_tb.v(104)
    output _cvpt_2274;   // oc8051_tb.v(104)
    output _cvpt_2275;   // oc8051_tb.v(104)
    output _cvpt_2276;   // oc8051_tb.v(104)
    output _cvpt_2277;   // oc8051_tb.v(104)
    output _cvpt_2278;   // oc8051_tb.v(104)
    output _cvpt_2279;   // oc8051_tb.v(104)
    output _cvpt_2280;   // oc8051_tb.v(104)
    output _cvpt_2281;   // oc8051_tb.v(104)
    output _cvpt_2282;   // oc8051_tb.v(104)
    output _cvpt_2283;   // oc8051_tb.v(104)
    output _cvpt_2284;   // oc8051_tb.v(104)
    output _cvpt_2285;   // oc8051_tb.v(104)
    output _cvpt_2286;   // oc8051_tb.v(104)
    output _cvpt_2287;   // oc8051_tb.v(104)
    output _cvpt_2288;   // oc8051_tb.v(104)
    output _cvpt_2289;   // oc8051_tb.v(104)
    output _cvpt_2290;   // oc8051_tb.v(104)
    output _cvpt_2291;   // oc8051_tb.v(104)
    output _cvpt_2292;   // oc8051_tb.v(104)
    output _cvpt_2293;   // oc8051_tb.v(104)
    output _cvpt_2294;   // oc8051_tb.v(104)
    output _cvpt_2295;   // oc8051_tb.v(104)
    output _cvpt_2296;   // oc8051_tb.v(104)
    output _cvpt_2297;   // oc8051_tb.v(104)
    output _cvpt_2298;   // oc8051_tb.v(104)
    output _cvpt_2299;   // oc8051_tb.v(104)
    output _cvpt_2300;   // oc8051_tb.v(104)
    output _cvpt_2301;   // oc8051_tb.v(104)
    output _cvpt_2302;   // oc8051_tb.v(104)
    output _cvpt_2303;   // oc8051_tb.v(104)
    output _cvpt_2304;   // oc8051_tb.v(104)
    output _cvpt_2305;   // oc8051_tb.v(104)
    output _cvpt_2306;   // oc8051_tb.v(104)
    output _cvpt_2307;   // oc8051_tb.v(104)
    output _cvpt_2308;   // oc8051_tb.v(104)
    output _cvpt_2309;   // oc8051_tb.v(104)
    output _cvpt_2310;   // oc8051_tb.v(104)
    output _cvpt_2311;   // oc8051_tb.v(104)
    output _cvpt_2312;   // oc8051_tb.v(104)
    output _cvpt_2313;   // oc8051_tb.v(104)
    output _cvpt_2314;   // oc8051_tb.v(104)
    output _cvpt_2315;   // oc8051_tb.v(104)
    output _cvpt_2316;   // oc8051_tb.v(104)
    output _cvpt_2317;   // oc8051_tb.v(104)
    output _cvpt_2318;   // oc8051_tb.v(104)
    output _cvpt_2319;   // oc8051_tb.v(104)
    output _cvpt_2320;   // oc8051_tb.v(104)
    output _cvpt_2321;   // oc8051_tb.v(104)
    output _cvpt_2322;   // oc8051_tb.v(104)
    output _cvpt_2323;   // oc8051_tb.v(104)
    output _cvpt_2324;   // oc8051_tb.v(104)
    output _cvpt_2325;   // oc8051_tb.v(104)
    output _cvpt_2326;   // oc8051_tb.v(104)
    output _cvpt_2327;   // oc8051_tb.v(104)
    output _cvpt_2328;   // oc8051_tb.v(104)
    output _cvpt_2329;   // oc8051_tb.v(104)
    output _cvpt_2330;   // oc8051_tb.v(104)
    output _cvpt_2331;   // oc8051_tb.v(104)
    output _cvpt_2332;   // oc8051_tb.v(104)
    output _cvpt_2333;   // oc8051_tb.v(104)
    output _cvpt_2334;   // oc8051_tb.v(104)
    output _cvpt_2335;   // oc8051_tb.v(104)
    output _cvpt_2336;   // oc8051_tb.v(104)
    output _cvpt_2337;   // oc8051_tb.v(104)
    output _cvpt_2338;   // oc8051_tb.v(104)
    output _cvpt_2339;   // oc8051_tb.v(104)
    output _cvpt_2340;   // oc8051_tb.v(104)
    output _cvpt_2341;   // oc8051_tb.v(104)
    output _cvpt_2342;   // oc8051_tb.v(104)
    output _cvpt_2343;   // oc8051_tb.v(104)
    output _cvpt_2344;   // oc8051_tb.v(104)
    output _cvpt_2345;   // oc8051_tb.v(104)
    output _cvpt_2346;   // oc8051_tb.v(104)
    output _cvpt_2347;   // oc8051_tb.v(104)
    output _cvpt_2348;   // oc8051_tb.v(104)
    output _cvpt_2349;   // oc8051_tb.v(104)
    output _cvpt_2350;   // oc8051_tb.v(104)
    output _cvpt_2351;   // oc8051_tb.v(104)
    output _cvpt_2352;   // oc8051_tb.v(104)
    output _cvpt_2353;   // oc8051_tb.v(104)
    output _cvpt_2354;   // oc8051_tb.v(104)
    output _cvpt_2355;   // oc8051_tb.v(104)
    output _cvpt_2356;   // oc8051_tb.v(104)
    output _cvpt_2357;   // oc8051_tb.v(104)
    output _cvpt_2358;   // oc8051_tb.v(104)
    output _cvpt_2359;   // oc8051_tb.v(104)
    output _cvpt_2360;   // oc8051_tb.v(104)
    output _cvpt_2361;   // oc8051_tb.v(104)
    output _cvpt_2362;   // oc8051_tb.v(104)
    output _cvpt_2363;   // oc8051_tb.v(104)
    output _cvpt_2364;   // oc8051_tb.v(104)
    output _cvpt_2365;   // oc8051_tb.v(104)
    output _cvpt_2366;   // oc8051_tb.v(104)
    output _cvpt_2367;   // oc8051_tb.v(104)
    output _cvpt_2368;   // oc8051_tb.v(104)
    output _cvpt_2369;   // oc8051_tb.v(104)
    output _cvpt_2370;   // oc8051_tb.v(104)
    output _cvpt_2371;   // oc8051_tb.v(104)
    output _cvpt_2372;   // oc8051_tb.v(104)
    output _cvpt_2373;   // oc8051_tb.v(104)
    output _cvpt_2374;   // oc8051_tb.v(104)
    output _cvpt_2375;   // oc8051_tb.v(104)
    output _cvpt_2376;   // oc8051_tb.v(104)
    output _cvpt_2377;   // oc8051_tb.v(104)
    output _cvpt_2378;   // oc8051_tb.v(104)
    output _cvpt_2379;   // oc8051_tb.v(104)
    output _cvpt_2380;   // oc8051_tb.v(104)
    output _cvpt_2381;   // oc8051_tb.v(104)
    output _cvpt_2382;   // oc8051_tb.v(104)
    output _cvpt_2383;   // oc8051_tb.v(104)
    output _cvpt_2384;   // oc8051_tb.v(104)
    output _cvpt_2385;   // oc8051_tb.v(104)
    output _cvpt_2386;   // oc8051_tb.v(104)
    output _cvpt_2387;   // oc8051_tb.v(104)
    output _cvpt_2388;   // oc8051_tb.v(104)
    output _cvpt_2389;   // oc8051_tb.v(104)
    output _cvpt_2390;   // oc8051_tb.v(104)
    output _cvpt_2391;   // oc8051_tb.v(104)
    output _cvpt_2392;   // oc8051_tb.v(104)
    output _cvpt_2393;   // oc8051_tb.v(104)
    output _cvpt_2394;   // oc8051_tb.v(104)
    output _cvpt_2395;   // oc8051_tb.v(104)
    output _cvpt_2396;   // oc8051_tb.v(104)
    output _cvpt_2397;   // oc8051_tb.v(104)
    output _cvpt_2398;   // oc8051_tb.v(104)
    output _cvpt_2399;   // oc8051_tb.v(104)
    output _cvpt_2400;   // oc8051_tb.v(104)
    output _cvpt_2401;   // oc8051_tb.v(104)
    output _cvpt_2402;   // oc8051_tb.v(104)
    output _cvpt_2403;   // oc8051_tb.v(104)
    output _cvpt_2404;   // oc8051_tb.v(104)
    output _cvpt_2405;   // oc8051_tb.v(104)
    output _cvpt_2406;   // oc8051_tb.v(104)
    output _cvpt_2407;   // oc8051_tb.v(104)
    output _cvpt_2408;   // oc8051_tb.v(104)
    output _cvpt_2409;   // oc8051_tb.v(104)
    output _cvpt_2410;   // oc8051_tb.v(104)
    output _cvpt_2411;   // oc8051_tb.v(104)
    output _cvpt_2412;   // oc8051_tb.v(104)
    output _cvpt_2413;   // oc8051_tb.v(104)
    output _cvpt_2414;   // oc8051_tb.v(104)
    output _cvpt_2415;   // oc8051_tb.v(104)
    output _cvpt_2416;   // oc8051_tb.v(104)
    output _cvpt_2417;   // oc8051_tb.v(104)
    output _cvpt_2418;   // oc8051_tb.v(104)
    output _cvpt_2419;   // oc8051_tb.v(104)
    output _cvpt_2420;   // oc8051_tb.v(104)
    output _cvpt_2421;   // oc8051_tb.v(104)
    output _cvpt_2422;   // oc8051_tb.v(104)
    output _cvpt_2423;   // oc8051_tb.v(104)
    output _cvpt_2424;   // oc8051_tb.v(104)
    output _cvpt_2425;   // oc8051_tb.v(104)
    output _cvpt_2426;   // oc8051_tb.v(104)
    output _cvpt_2427;   // oc8051_tb.v(104)
    output _cvpt_2428;   // oc8051_tb.v(104)
    output _cvpt_2429;   // oc8051_tb.v(104)
    output _cvpt_2430;   // oc8051_tb.v(104)
    output _cvpt_2431;   // oc8051_tb.v(104)
    output _cvpt_2432;   // oc8051_tb.v(104)
    output _cvpt_2433;   // oc8051_tb.v(104)
    output _cvpt_2434;   // oc8051_tb.v(104)
    output _cvpt_2435;   // oc8051_tb.v(104)
    output _cvpt_2436;   // oc8051_tb.v(104)
    output _cvpt_2437;   // oc8051_tb.v(104)
    output _cvpt_2438;   // oc8051_tb.v(104)
    output _cvpt_2439;   // oc8051_tb.v(104)
    output _cvpt_2440;   // oc8051_tb.v(104)
    output _cvpt_2441;   // oc8051_tb.v(104)
    output _cvpt_2442;   // oc8051_tb.v(104)
    output _cvpt_2443;   // oc8051_tb.v(104)
    output _cvpt_2444;   // oc8051_tb.v(104)
    output _cvpt_2445;   // oc8051_tb.v(104)
    output _cvpt_2446;   // oc8051_tb.v(104)
    output _cvpt_2447;   // oc8051_tb.v(104)
    output _cvpt_2448;   // oc8051_tb.v(104)
    output _cvpt_2449;   // oc8051_tb.v(104)
    output _cvpt_2450;   // oc8051_tb.v(104)
    output _cvpt_2451;   // oc8051_tb.v(104)
    output _cvpt_2452;   // oc8051_tb.v(104)
    output _cvpt_2453;   // oc8051_tb.v(104)
    output _cvpt_2454;   // oc8051_tb.v(104)
    output _cvpt_2455;   // oc8051_tb.v(104)
    output _cvpt_2456;   // oc8051_tb.v(104)
    output _cvpt_2457;   // oc8051_tb.v(104)
    output _cvpt_2458;   // oc8051_tb.v(104)
    output _cvpt_2459;   // oc8051_tb.v(104)
    output _cvpt_2460;   // oc8051_tb.v(104)
    output _cvpt_2461;   // oc8051_tb.v(104)
    output _cvpt_2462;   // oc8051_tb.v(104)
    output _cvpt_2463;   // oc8051_tb.v(104)
    output _cvpt_2464;   // oc8051_tb.v(104)
    output _cvpt_2465;   // oc8051_tb.v(104)
    output _cvpt_2466;   // oc8051_tb.v(104)
    output _cvpt_2467;   // oc8051_tb.v(104)
    output _cvpt_2468;   // oc8051_tb.v(104)
    output _cvpt_2469;   // oc8051_tb.v(104)
    output _cvpt_2470;   // oc8051_tb.v(104)
    output _cvpt_2471;   // oc8051_tb.v(104)
    output _cvpt_2472;   // oc8051_tb.v(104)
    output _cvpt_2473;   // oc8051_tb.v(104)
    output _cvpt_2474;   // oc8051_tb.v(104)
    output _cvpt_2475;   // oc8051_tb.v(104)
    output _cvpt_2476;   // oc8051_tb.v(104)
    output _cvpt_2477;   // oc8051_tb.v(104)
    output _cvpt_2478;   // oc8051_tb.v(104)
    output _cvpt_2479;   // oc8051_tb.v(104)
    output _cvpt_2480;   // oc8051_tb.v(104)
    output _cvpt_2481;   // oc8051_tb.v(104)
    output _cvpt_2482;   // oc8051_tb.v(104)
    output _cvpt_2483;   // oc8051_tb.v(104)
    output _cvpt_2484;   // oc8051_tb.v(104)
    output _cvpt_2485;   // oc8051_tb.v(104)
    output _cvpt_2486;   // oc8051_tb.v(104)
    output _cvpt_2487;   // oc8051_tb.v(104)
    output _cvpt_2488;   // oc8051_tb.v(104)
    output _cvpt_2489;   // oc8051_tb.v(104)
    output _cvpt_2490;   // oc8051_tb.v(104)
    output _cvpt_2491;   // oc8051_tb.v(104)
    output _cvpt_2492;   // oc8051_tb.v(104)
    output _cvpt_2493;   // oc8051_tb.v(104)
    output _cvpt_2494;   // oc8051_tb.v(104)
    output _cvpt_2495;   // oc8051_tb.v(104)
    output _cvpt_2496;   // oc8051_tb.v(104)
    output _cvpt_2497;   // oc8051_tb.v(104)
    output _cvpt_2498;   // oc8051_tb.v(104)
    output _cvpt_2499;   // oc8051_tb.v(104)
    output _cvpt_2500;   // oc8051_tb.v(104)
    output _cvpt_2501;   // oc8051_tb.v(104)
    output _cvpt_2502;   // oc8051_tb.v(104)
    output _cvpt_2503;   // oc8051_tb.v(104)
    output _cvpt_2504;   // oc8051_tb.v(104)
    output _cvpt_2505;   // oc8051_tb.v(104)
    output _cvpt_2506;   // oc8051_tb.v(104)
    output _cvpt_2507;   // oc8051_tb.v(104)
    output _cvpt_2508;   // oc8051_tb.v(104)
    output _cvpt_2509;   // oc8051_tb.v(104)
    output _cvpt_2510;   // oc8051_tb.v(104)
    output _cvpt_2511;   // oc8051_tb.v(104)
    output _cvpt_2512;   // oc8051_tb.v(104)
    output _cvpt_2513;   // oc8051_tb.v(104)
    output _cvpt_2514;   // oc8051_tb.v(104)
    output _cvpt_2515;   // oc8051_tb.v(104)
    output _cvpt_2516;   // oc8051_tb.v(104)
    output _cvpt_2517;   // oc8051_tb.v(104)
    output _cvpt_2518;   // oc8051_tb.v(104)
    output _cvpt_2519;   // oc8051_tb.v(104)
    output _cvpt_2520;   // oc8051_tb.v(104)
    output _cvpt_2521;   // oc8051_tb.v(104)
    output _cvpt_2522;   // oc8051_tb.v(104)
    output _cvpt_2523;   // oc8051_tb.v(104)
    output _cvpt_2524;   // oc8051_tb.v(104)
    output _cvpt_2525;   // oc8051_tb.v(104)
    output _cvpt_2526;   // oc8051_tb.v(104)
    output _cvpt_2527;   // oc8051_tb.v(104)
    output _cvpt_2528;   // oc8051_tb.v(104)
    output _cvpt_2529;   // oc8051_tb.v(104)
    output _cvpt_2530;   // oc8051_tb.v(104)
    output _cvpt_2531;   // oc8051_tb.v(104)
    output _cvpt_2532;   // oc8051_tb.v(104)
    output _cvpt_2533;   // oc8051_tb.v(104)
    output _cvpt_2534;   // oc8051_tb.v(104)
    output _cvpt_2535;   // oc8051_tb.v(104)
    output _cvpt_2536;   // oc8051_tb.v(104)
    output _cvpt_2537;   // oc8051_tb.v(104)
    output _cvpt_2538;   // oc8051_tb.v(104)
    output _cvpt_2539;   // oc8051_tb.v(104)
    output _cvpt_2540;   // oc8051_tb.v(104)
    output _cvpt_2541;   // oc8051_tb.v(104)
    output _cvpt_2542;   // oc8051_tb.v(104)
    output _cvpt_2543;   // oc8051_tb.v(104)
    output _cvpt_2544;   // oc8051_tb.v(104)
    output _cvpt_2545;   // oc8051_tb.v(104)
    output _cvpt_2546;   // oc8051_tb.v(104)
    output _cvpt_2547;   // oc8051_tb.v(104)
    output _cvpt_2548;   // oc8051_tb.v(104)
    output _cvpt_2549;   // oc8051_tb.v(104)
    output _cvpt_2550;   // oc8051_tb.v(104)
    output _cvpt_2551;   // oc8051_tb.v(104)
    output _cvpt_2552;   // oc8051_tb.v(104)
    output _cvpt_2553;   // oc8051_tb.v(104)
    output _cvpt_2554;   // oc8051_tb.v(104)
    output _cvpt_2555;   // oc8051_tb.v(104)
    output _cvpt_2556;   // oc8051_tb.v(104)
    output _cvpt_2557;   // oc8051_tb.v(104)
    output _cvpt_2558;   // oc8051_tb.v(104)
    output _cvpt_2559;   // oc8051_tb.v(104)
    output _cvpt_2560;   // oc8051_tb.v(104)
    output _cvpt_2561;   // oc8051_tb.v(104)
    output _cvpt_2562;   // oc8051_tb.v(104)
    output _cvpt_2563;   // oc8051_tb.v(104)
    output _cvpt_2564;   // oc8051_tb.v(104)
    output _cvpt_2565;   // oc8051_tb.v(104)
    output _cvpt_2566;   // oc8051_tb.v(104)
    output _cvpt_2567;   // oc8051_tb.v(104)
    output _cvpt_2568;   // oc8051_tb.v(104)
    output _cvpt_2569;   // oc8051_tb.v(104)
    output _cvpt_2570;   // oc8051_tb.v(104)
    output _cvpt_2571;   // oc8051_tb.v(104)
    output _cvpt_2572;   // oc8051_tb.v(104)
    output _cvpt_2573;   // oc8051_tb.v(104)
    output _cvpt_2574;   // oc8051_tb.v(104)
    output _cvpt_2575;   // oc8051_tb.v(104)
    output _cvpt_2576;   // oc8051_tb.v(104)
    output _cvpt_2577;   // oc8051_tb.v(104)
    output _cvpt_2578;   // oc8051_tb.v(104)
    output _cvpt_2579;   // oc8051_tb.v(104)
    output _cvpt_2580;   // oc8051_tb.v(104)
    output _cvpt_2581;   // oc8051_tb.v(104)
    output _cvpt_2582;   // oc8051_tb.v(104)
    output _cvpt_2583;   // oc8051_tb.v(104)
    output _cvpt_2584;   // oc8051_tb.v(104)
    output _cvpt_2585;   // oc8051_tb.v(104)
    output _cvpt_2586;   // oc8051_tb.v(104)
    output _cvpt_2587;   // oc8051_tb.v(104)
    output _cvpt_2588;   // oc8051_tb.v(104)
    output _cvpt_2589;   // oc8051_tb.v(104)
    output _cvpt_2590;   // oc8051_tb.v(104)
    output _cvpt_2591;   // oc8051_tb.v(104)
    output _cvpt_2592;   // oc8051_tb.v(104)
    output _cvpt_2593;   // oc8051_tb.v(104)
    output _cvpt_2594;   // oc8051_tb.v(104)
    output _cvpt_2595;   // oc8051_tb.v(104)
    output _cvpt_2596;   // oc8051_tb.v(104)
    output _cvpt_2597;   // oc8051_tb.v(104)
    output _cvpt_2598;   // oc8051_tb.v(104)
    output _cvpt_2599;   // oc8051_tb.v(104)
    output _cvpt_2600;   // oc8051_tb.v(104)
    output _cvpt_2601;   // oc8051_tb.v(104)
    output _cvpt_2602;   // oc8051_tb.v(104)
    output _cvpt_2603;   // oc8051_tb.v(104)
    output _cvpt_2604;   // oc8051_tb.v(104)
    output _cvpt_2605;   // oc8051_tb.v(104)
    output _cvpt_2606;   // oc8051_tb.v(104)
    output _cvpt_2607;   // oc8051_tb.v(104)
    output _cvpt_2608;   // oc8051_tb.v(104)
    output _cvpt_2609;   // oc8051_tb.v(104)
    output _cvpt_2610;   // oc8051_tb.v(104)
    output _cvpt_2611;   // oc8051_tb.v(104)
    output _cvpt_2612;   // oc8051_tb.v(104)
    output _cvpt_2613;   // oc8051_tb.v(104)
    output _cvpt_2614;   // oc8051_tb.v(104)
    output _cvpt_2615;   // oc8051_tb.v(104)
    output _cvpt_2616;   // oc8051_tb.v(104)
    output _cvpt_2617;   // oc8051_tb.v(104)
    output _cvpt_2618;   // oc8051_tb.v(104)
    output _cvpt_2619;   // oc8051_tb.v(104)
    output _cvpt_2620;   // oc8051_tb.v(104)
    output _cvpt_2621;   // oc8051_tb.v(104)
    output _cvpt_2622;   // oc8051_tb.v(104)
    output _cvpt_2623;   // oc8051_tb.v(104)
    output _cvpt_2624;   // oc8051_tb.v(104)
    output _cvpt_2625;   // oc8051_tb.v(104)
    output _cvpt_2626;   // oc8051_tb.v(104)
    output _cvpt_2627;   // oc8051_tb.v(104)
    output _cvpt_2628;   // oc8051_tb.v(104)
    output _cvpt_2629;   // oc8051_tb.v(104)
    output _cvpt_2630;   // oc8051_tb.v(104)
    output _cvpt_2631;   // oc8051_tb.v(104)
    output _cvpt_2632;   // oc8051_tb.v(104)
    output _cvpt_2633;   // oc8051_tb.v(104)
    output _cvpt_2634;   // oc8051_tb.v(104)
    output _cvpt_2635;   // oc8051_tb.v(104)
    output _cvpt_2636;   // oc8051_tb.v(104)
    output _cvpt_2637;   // oc8051_tb.v(104)
    output _cvpt_2638;   // oc8051_tb.v(104)
    output _cvpt_2639;   // oc8051_tb.v(104)
    output _cvpt_2640;   // oc8051_tb.v(104)
    output _cvpt_2641;   // oc8051_tb.v(104)
    output _cvpt_2642;   // oc8051_tb.v(104)
    output _cvpt_2643;   // oc8051_tb.v(104)
    output _cvpt_2644;   // oc8051_tb.v(104)
    output _cvpt_2645;   // oc8051_tb.v(104)
    output _cvpt_2646;   // oc8051_tb.v(104)
    output _cvpt_2647;   // oc8051_tb.v(104)
    output _cvpt_2648;   // oc8051_tb.v(104)
    output _cvpt_2649;   // oc8051_tb.v(104)
    output _cvpt_2650;   // oc8051_tb.v(104)
    output _cvpt_2651;   // oc8051_tb.v(104)
    output _cvpt_2652;   // oc8051_tb.v(104)
    output _cvpt_2653;   // oc8051_tb.v(104)
    output _cvpt_2654;   // oc8051_tb.v(104)
    output _cvpt_2655;   // oc8051_tb.v(104)
    output _cvpt_2656;   // oc8051_tb.v(104)
    output _cvpt_2657;   // oc8051_tb.v(104)
    output _cvpt_2658;   // oc8051_tb.v(104)
    output _cvpt_2659;   // oc8051_tb.v(104)
    output _cvpt_2660;   // oc8051_tb.v(104)
    output _cvpt_2661;   // oc8051_tb.v(104)
    output _cvpt_2662;   // oc8051_tb.v(104)
    output _cvpt_2663;   // oc8051_tb.v(104)
    output _cvpt_2664;   // oc8051_tb.v(104)
    output _cvpt_2665;   // oc8051_tb.v(104)
    output _cvpt_2666;   // oc8051_tb.v(104)
    output _cvpt_2667;   // oc8051_tb.v(104)
    output _cvpt_2668;   // oc8051_tb.v(104)
    output _cvpt_2669;   // oc8051_tb.v(104)
    output _cvpt_2670;   // oc8051_tb.v(104)
    output _cvpt_2671;   // oc8051_tb.v(104)
    output _cvpt_2672;   // oc8051_tb.v(104)
    output _cvpt_2673;   // oc8051_tb.v(104)
    output _cvpt_2674;   // oc8051_tb.v(104)
    output _cvpt_2675;   // oc8051_tb.v(104)
    output _cvpt_2676;   // oc8051_tb.v(104)
    output _cvpt_2677;   // oc8051_tb.v(104)
    output _cvpt_2678;   // oc8051_tb.v(104)
    output _cvpt_2679;   // oc8051_tb.v(104)
    output _cvpt_2680;   // oc8051_tb.v(104)
    output _cvpt_2681;   // oc8051_tb.v(104)
    output _cvpt_2682;   // oc8051_tb.v(104)
    output _cvpt_2683;   // oc8051_tb.v(104)
    output _cvpt_2684;   // oc8051_tb.v(104)
    output _cvpt_2685;   // oc8051_tb.v(104)
    output _cvpt_2686;   // oc8051_tb.v(104)
    output _cvpt_2687;   // oc8051_tb.v(104)
    output _cvpt_2688;   // oc8051_tb.v(104)
    output _cvpt_2689;   // oc8051_tb.v(104)
    output _cvpt_2690;   // oc8051_tb.v(104)
    output _cvpt_2691;   // oc8051_tb.v(104)
    output _cvpt_2692;   // oc8051_tb.v(104)
    output _cvpt_2693;   // oc8051_tb.v(104)
    output _cvpt_2694;   // oc8051_tb.v(104)
    output _cvpt_2695;   // oc8051_tb.v(104)
    output _cvpt_2696;   // oc8051_tb.v(104)
    output _cvpt_2697;   // oc8051_tb.v(104)
    output _cvpt_2698;   // oc8051_tb.v(104)
    output _cvpt_2699;   // oc8051_tb.v(104)
    output _cvpt_2700;   // oc8051_tb.v(104)
    output _cvpt_2701;   // oc8051_tb.v(104)
    output _cvpt_2702;   // oc8051_tb.v(104)
    output _cvpt_2703;   // oc8051_tb.v(104)
    output _cvpt_2704;   // oc8051_tb.v(104)
    output _cvpt_2705;   // oc8051_tb.v(104)
    output _cvpt_2706;   // oc8051_tb.v(104)
    output _cvpt_2707;   // oc8051_tb.v(104)
    output _cvpt_2708;   // oc8051_tb.v(104)
    output _cvpt_2709;   // oc8051_tb.v(104)
    output _cvpt_2710;   // oc8051_tb.v(104)
    output _cvpt_2711;   // oc8051_tb.v(104)
    output _cvpt_2712;   // oc8051_tb.v(104)
    output _cvpt_2713;   // oc8051_tb.v(104)
    output _cvpt_2714;   // oc8051_tb.v(104)
    output _cvpt_2715;   // oc8051_tb.v(104)
    output _cvpt_2716;   // oc8051_tb.v(104)
    output _cvpt_2717;   // oc8051_tb.v(104)
    output _cvpt_2718;   // oc8051_tb.v(104)
    output _cvpt_2719;   // oc8051_tb.v(104)
    output _cvpt_2720;   // oc8051_tb.v(104)
    output _cvpt_2721;   // oc8051_tb.v(104)
    output _cvpt_2722;   // oc8051_tb.v(104)
    output _cvpt_2723;   // oc8051_tb.v(104)
    output _cvpt_2724;   // oc8051_tb.v(104)
    output _cvpt_2725;   // oc8051_tb.v(104)
    output _cvpt_2726;   // oc8051_tb.v(104)
    output _cvpt_2727;   // oc8051_tb.v(104)
    output _cvpt_2728;   // oc8051_tb.v(104)
    output _cvpt_2729;   // oc8051_tb.v(104)
    output _cvpt_2730;   // oc8051_tb.v(104)
    output _cvpt_2731;   // oc8051_tb.v(104)
    output _cvpt_2732;   // oc8051_tb.v(104)
    output _cvpt_2733;   // oc8051_tb.v(104)
    output _cvpt_2734;   // oc8051_tb.v(104)
    output _cvpt_2735;   // oc8051_tb.v(104)
    output _cvpt_2736;   // oc8051_tb.v(104)
    output _cvpt_2737;   // oc8051_tb.v(104)
    output _cvpt_2738;   // oc8051_tb.v(104)
    output _cvpt_2739;   // oc8051_tb.v(104)
    output _cvpt_2740;   // oc8051_tb.v(104)
    output _cvpt_2741;   // oc8051_tb.v(104)
    output _cvpt_2742;   // oc8051_tb.v(104)
    output _cvpt_2743;   // oc8051_tb.v(104)
    output _cvpt_2744;   // oc8051_tb.v(104)
    output _cvpt_2745;   // oc8051_tb.v(104)
    output _cvpt_2746;   // oc8051_tb.v(104)
    output _cvpt_2747;   // oc8051_tb.v(104)
    output _cvpt_2748;   // oc8051_tb.v(104)
    output _cvpt_2749;   // oc8051_tb.v(104)
    output _cvpt_2750;   // oc8051_tb.v(104)
    output _cvpt_2751;   // oc8051_tb.v(104)
    output _cvpt_2752;   // oc8051_tb.v(104)
    output _cvpt_2753;   // oc8051_tb.v(104)
    output _cvpt_2754;   // oc8051_tb.v(104)
    output _cvpt_2755;   // oc8051_tb.v(104)
    output _cvpt_2756;   // oc8051_tb.v(104)
    output _cvpt_2757;   // oc8051_tb.v(104)
    output _cvpt_2758;   // oc8051_tb.v(104)
    output _cvpt_2759;   // oc8051_tb.v(104)
    output _cvpt_2760;   // oc8051_tb.v(104)
    output _cvpt_2761;   // oc8051_tb.v(104)
    output _cvpt_2762;   // oc8051_tb.v(104)
    output _cvpt_2763;   // oc8051_tb.v(104)
    output _cvpt_2764;   // oc8051_tb.v(104)
    output _cvpt_2765;   // oc8051_tb.v(104)
    output _cvpt_2766;   // oc8051_tb.v(104)
    output _cvpt_2767;   // oc8051_tb.v(104)
    output _cvpt_2768;   // oc8051_tb.v(104)
    output _cvpt_2769;   // oc8051_tb.v(104)
    output _cvpt_2770;   // oc8051_tb.v(104)
    output _cvpt_2771;   // oc8051_tb.v(104)
    output _cvpt_2772;   // oc8051_tb.v(104)
    output _cvpt_2773;   // oc8051_tb.v(104)
    output _cvpt_2774;   // oc8051_tb.v(104)
    output _cvpt_2775;   // oc8051_tb.v(104)
    output _cvpt_2776;   // oc8051_tb.v(104)
    output _cvpt_2777;   // oc8051_tb.v(104)
    output _cvpt_2778;   // oc8051_tb.v(104)
    output _cvpt_2779;   // oc8051_tb.v(104)
    output _cvpt_2780;   // oc8051_tb.v(104)
    output _cvpt_2781;   // oc8051_tb.v(104)
    output _cvpt_2782;   // oc8051_tb.v(104)
    output _cvpt_2783;   // oc8051_tb.v(104)
    output _cvpt_2784;   // oc8051_tb.v(104)
    output _cvpt_2785;   // oc8051_tb.v(104)
    output _cvpt_2786;   // oc8051_tb.v(104)
    output _cvpt_2787;   // oc8051_tb.v(104)
    output _cvpt_2788;   // oc8051_tb.v(104)
    output _cvpt_2789;   // oc8051_tb.v(104)
    output _cvpt_2790;   // oc8051_tb.v(104)
    output _cvpt_2791;   // oc8051_tb.v(104)
    output _cvpt_2792;   // oc8051_tb.v(104)
    output _cvpt_2793;   // oc8051_tb.v(104)
    output _cvpt_2794;   // oc8051_tb.v(104)
    output _cvpt_2795;   // oc8051_tb.v(104)
    output _cvpt_2796;   // oc8051_tb.v(104)
    output _cvpt_2797;   // oc8051_tb.v(104)
    output _cvpt_2798;   // oc8051_tb.v(104)
    output _cvpt_2799;   // oc8051_tb.v(104)
    output _cvpt_2800;   // oc8051_tb.v(104)
    output _cvpt_2801;   // oc8051_tb.v(104)
    output _cvpt_2802;   // oc8051_tb.v(104)
    output _cvpt_2803;   // oc8051_tb.v(104)
    output _cvpt_2804;   // oc8051_tb.v(104)
    output _cvpt_2805;   // oc8051_tb.v(104)
    output _cvpt_2806;   // oc8051_tb.v(104)
    output _cvpt_2807;   // oc8051_tb.v(104)
    output _cvpt_2808;   // oc8051_tb.v(104)
    output _cvpt_2809;   // oc8051_tb.v(104)
    output _cvpt_2810;   // oc8051_tb.v(104)
    output _cvpt_2811;   // oc8051_tb.v(104)
    output _cvpt_2812;   // oc8051_tb.v(104)
    output _cvpt_2813;   // oc8051_tb.v(104)
    output _cvpt_2814;   // oc8051_tb.v(104)
    output _cvpt_2815;   // oc8051_tb.v(104)
    output _cvpt_2816;   // oc8051_tb.v(104)
    output _cvpt_2817;   // oc8051_tb.v(104)
    output _cvpt_2818;   // oc8051_tb.v(104)
    output _cvpt_2819;   // oc8051_tb.v(104)
    output _cvpt_2820;   // oc8051_tb.v(104)
    output _cvpt_2821;   // oc8051_tb.v(104)
    output _cvpt_2822;   // oc8051_tb.v(104)
    output _cvpt_2823;   // oc8051_tb.v(104)
    output _cvpt_2824;   // oc8051_tb.v(104)
    output _cvpt_2825;   // oc8051_tb.v(104)
    output _cvpt_2826;   // oc8051_tb.v(104)
    output _cvpt_2827;   // oc8051_tb.v(104)
    output _cvpt_2828;   // oc8051_tb.v(104)
    output _cvpt_2829;   // oc8051_tb.v(104)
    output _cvpt_2830;   // oc8051_tb.v(104)
    output _cvpt_2831;   // oc8051_tb.v(104)
    output _cvpt_2832;   // oc8051_tb.v(104)
    output _cvpt_2833;   // oc8051_tb.v(104)
    output _cvpt_2834;   // oc8051_tb.v(104)
    output _cvpt_2835;   // oc8051_tb.v(104)
    output _cvpt_2836;   // oc8051_tb.v(104)
    output _cvpt_2837;   // oc8051_tb.v(104)
    output _cvpt_2838;   // oc8051_tb.v(104)
    output _cvpt_2839;   // oc8051_tb.v(104)
    output _cvpt_2840;   // oc8051_tb.v(104)
    output _cvpt_2841;   // oc8051_tb.v(104)
    output _cvpt_2842;   // oc8051_tb.v(104)
    output _cvpt_2843;   // oc8051_tb.v(104)
    output _cvpt_2844;   // oc8051_tb.v(104)
    output _cvpt_2845;   // oc8051_tb.v(104)
    output _cvpt_2846;   // oc8051_tb.v(104)
    output _cvpt_2847;   // oc8051_tb.v(104)
    output _cvpt_2848;   // oc8051_tb.v(104)
    output _cvpt_2849;   // oc8051_tb.v(104)
    output _cvpt_2850;   // oc8051_tb.v(104)
    output _cvpt_2851;   // oc8051_tb.v(104)
    output _cvpt_2852;   // oc8051_tb.v(104)
    output _cvpt_2853;   // oc8051_tb.v(104)
    output _cvpt_2854;   // oc8051_tb.v(104)
    output _cvpt_2855;   // oc8051_tb.v(104)
    output _cvpt_2856;   // oc8051_tb.v(104)
    output _cvpt_2857;   // oc8051_tb.v(104)
    output _cvpt_2858;   // oc8051_tb.v(104)
    output _cvpt_2859;   // oc8051_tb.v(104)
    output _cvpt_2860;   // oc8051_tb.v(104)
    output _cvpt_2861;   // oc8051_tb.v(104)
    output _cvpt_2862;   // oc8051_tb.v(104)
    output _cvpt_2863;   // oc8051_tb.v(104)
    output _cvpt_2864;   // oc8051_tb.v(104)
    output _cvpt_2865;   // oc8051_tb.v(104)
    output _cvpt_2866;   // oc8051_tb.v(104)
    output _cvpt_2867;   // oc8051_tb.v(104)
    output _cvpt_2868;   // oc8051_tb.v(104)
    output _cvpt_2869;   // oc8051_tb.v(104)
    output _cvpt_2870;   // oc8051_tb.v(104)
    output _cvpt_2871;   // oc8051_tb.v(104)
    output _cvpt_2872;   // oc8051_tb.v(104)
    output _cvpt_2873;   // oc8051_tb.v(104)
    output _cvpt_2874;   // oc8051_tb.v(104)
    output _cvpt_2875;   // oc8051_tb.v(104)
    output _cvpt_2876;   // oc8051_tb.v(104)
    output _cvpt_2877;   // oc8051_tb.v(104)
    output _cvpt_2878;   // oc8051_tb.v(104)
    output _cvpt_2879;   // oc8051_tb.v(104)
    output _cvpt_2880;   // oc8051_tb.v(104)
    output _cvpt_2881;   // oc8051_tb.v(104)
    output _cvpt_2882;   // oc8051_tb.v(104)
    output _cvpt_2883;   // oc8051_tb.v(104)
    output _cvpt_2884;   // oc8051_tb.v(104)
    output _cvpt_2885;   // oc8051_tb.v(104)
    output _cvpt_2886;   // oc8051_tb.v(104)
    output _cvpt_2887;   // oc8051_tb.v(104)
    output _cvpt_2888;   // oc8051_tb.v(104)
    output _cvpt_2889;   // oc8051_tb.v(104)
    output _cvpt_2890;   // oc8051_tb.v(104)
    output _cvpt_2891;   // oc8051_tb.v(104)
    output _cvpt_2892;   // oc8051_tb.v(104)
    output _cvpt_2893;   // oc8051_tb.v(104)
    output _cvpt_2894;   // oc8051_tb.v(104)
    output _cvpt_2895;   // oc8051_tb.v(104)
    output _cvpt_2896;   // oc8051_tb.v(104)
    output _cvpt_2897;   // oc8051_tb.v(104)
    output _cvpt_2898;   // oc8051_tb.v(104)
    output _cvpt_2899;   // oc8051_tb.v(104)
    output _cvpt_2900;   // oc8051_tb.v(104)
    output _cvpt_2901;   // oc8051_tb.v(104)
    output _cvpt_2902;   // oc8051_tb.v(104)
    output _cvpt_2903;   // oc8051_tb.v(104)
    output _cvpt_2904;   // oc8051_tb.v(104)
    output _cvpt_2905;   // oc8051_tb.v(104)
    output _cvpt_2906;   // oc8051_tb.v(104)
    output _cvpt_2907;   // oc8051_tb.v(104)
    output _cvpt_2908;   // oc8051_tb.v(104)
    output _cvpt_2909;   // oc8051_tb.v(104)
    output _cvpt_2910;   // oc8051_tb.v(104)
    output _cvpt_2911;   // oc8051_tb.v(104)
    output _cvpt_2912;   // oc8051_tb.v(104)
    output _cvpt_2913;   // oc8051_tb.v(104)
    output _cvpt_2914;   // oc8051_tb.v(104)
    output _cvpt_2915;   // oc8051_tb.v(104)
    output _cvpt_2916;   // oc8051_tb.v(104)
    output _cvpt_2917;   // oc8051_tb.v(104)
    output _cvpt_2918;   // oc8051_tb.v(104)
    output _cvpt_2919;   // oc8051_tb.v(104)
    output _cvpt_2920;   // oc8051_tb.v(104)
    output _cvpt_2921;   // oc8051_tb.v(104)
    output _cvpt_2922;   // oc8051_tb.v(104)
    output _cvpt_2923;   // oc8051_tb.v(104)
    output _cvpt_2924;   // oc8051_tb.v(104)
    output _cvpt_2925;   // oc8051_tb.v(104)
    output _cvpt_2926;   // oc8051_tb.v(104)
    output _cvpt_2927;   // oc8051_tb.v(104)
    output _cvpt_2928;   // oc8051_tb.v(104)
    output _cvpt_2929;   // oc8051_tb.v(104)
    output _cvpt_2930;   // oc8051_tb.v(104)
    output _cvpt_2931;   // oc8051_tb.v(104)
    output _cvpt_2932;   // oc8051_tb.v(104)
    output _cvpt_2933;   // oc8051_tb.v(104)
    output _cvpt_2934;   // oc8051_tb.v(104)
    output _cvpt_2935;   // oc8051_tb.v(104)
    output _cvpt_2936;   // oc8051_tb.v(104)
    output _cvpt_2937;   // oc8051_tb.v(104)
    output _cvpt_2938;   // oc8051_tb.v(104)
    output _cvpt_2939;   // oc8051_tb.v(104)
    output _cvpt_2940;   // oc8051_tb.v(104)
    output _cvpt_2941;   // oc8051_tb.v(104)
    output _cvpt_2942;   // oc8051_tb.v(104)
    output _cvpt_2943;   // oc8051_tb.v(104)
    output _cvpt_2944;   // oc8051_tb.v(104)
    output _cvpt_2945;   // oc8051_tb.v(104)
    output _cvpt_2946;   // oc8051_tb.v(104)
    output _cvpt_2947;   // oc8051_tb.v(104)
    output _cvpt_2948;   // oc8051_tb.v(104)
    output _cvpt_2949;   // oc8051_tb.v(104)
    output _cvpt_2950;   // oc8051_tb.v(104)
    output _cvpt_2951;   // oc8051_tb.v(104)
    output _cvpt_2952;   // oc8051_tb.v(104)
    output _cvpt_2953;   // oc8051_tb.v(104)
    output _cvpt_2954;   // oc8051_tb.v(104)
    output _cvpt_2955;   // oc8051_tb.v(104)
    output _cvpt_2956;   // oc8051_tb.v(104)
    output _cvpt_2957;   // oc8051_tb.v(104)
    output _cvpt_2958;   // oc8051_tb.v(104)
    output _cvpt_2959;   // oc8051_tb.v(104)
    output _cvpt_2960;   // oc8051_tb.v(104)
    output _cvpt_2961;   // oc8051_tb.v(104)
    output _cvpt_2962;   // oc8051_tb.v(104)
    output _cvpt_2963;   // oc8051_tb.v(104)
    output _cvpt_2964;   // oc8051_tb.v(104)
    output _cvpt_2965;   // oc8051_tb.v(104)
    output _cvpt_2966;   // oc8051_tb.v(104)
    output _cvpt_2967;   // oc8051_tb.v(104)
    output _cvpt_2968;   // oc8051_tb.v(104)
    output _cvpt_2969;   // oc8051_tb.v(104)
    output _cvpt_2970;   // oc8051_tb.v(104)
    output _cvpt_2971;   // oc8051_tb.v(104)
    output _cvpt_2972;   // oc8051_tb.v(104)
    output _cvpt_2973;   // oc8051_tb.v(104)
    output _cvpt_2974;   // oc8051_tb.v(104)
    output _cvpt_2975;   // oc8051_tb.v(104)
    output _cvpt_2976;   // oc8051_tb.v(104)
    output _cvpt_2977;   // oc8051_tb.v(104)
    output _cvpt_2978;   // oc8051_tb.v(104)
    output _cvpt_2979;   // oc8051_tb.v(104)
    output _cvpt_2980;   // oc8051_tb.v(104)
    output _cvpt_2981;   // oc8051_tb.v(104)
    output _cvpt_2982;   // oc8051_tb.v(104)
    output _cvpt_2983;   // oc8051_tb.v(104)
    output _cvpt_2984;   // oc8051_tb.v(104)
    output _cvpt_2985;   // oc8051_tb.v(104)
    output _cvpt_2986;   // oc8051_tb.v(104)
    output _cvpt_2987;   // oc8051_tb.v(104)
    output _cvpt_2988;   // oc8051_tb.v(104)
    output _cvpt_2989;   // oc8051_tb.v(104)
    output _cvpt_2990;   // oc8051_tb.v(104)
    output _cvpt_2991;   // oc8051_tb.v(104)
    output _cvpt_2992;   // oc8051_tb.v(104)
    output _cvpt_2993;   // oc8051_tb.v(104)
    output _cvpt_2994;   // oc8051_tb.v(104)
    output _cvpt_2995;   // oc8051_tb.v(104)
    output _cvpt_2996;   // oc8051_tb.v(104)
    output _cvpt_2997;   // oc8051_tb.v(104)
    output _cvpt_2998;   // oc8051_tb.v(104)
    output _cvpt_2999;   // oc8051_tb.v(104)
    output _cvpt_3000;   // oc8051_tb.v(104)
    output _cvpt_3001;   // oc8051_tb.v(104)
    output _cvpt_3002;   // oc8051_tb.v(104)
    output _cvpt_3003;   // oc8051_tb.v(104)
    output _cvpt_3004;   // oc8051_tb.v(104)
    output _cvpt_3005;   // oc8051_tb.v(104)
    output _cvpt_3006;   // oc8051_tb.v(104)
    output _cvpt_3007;   // oc8051_tb.v(104)
    output _cvpt_3008;   // oc8051_tb.v(104)
    output _cvpt_3009;   // oc8051_tb.v(104)
    output _cvpt_3010;   // oc8051_tb.v(104)
    output _cvpt_3011;   // oc8051_tb.v(104)
    output _cvpt_3012;   // oc8051_tb.v(104)
    output _cvpt_3013;   // oc8051_tb.v(104)
    output _cvpt_3014;   // oc8051_tb.v(104)
    output _cvpt_3015;   // oc8051_tb.v(104)
    output _cvpt_3016;   // oc8051_tb.v(104)
    output _cvpt_3017;   // oc8051_tb.v(104)
    output _cvpt_3018;   // oc8051_tb.v(104)
    output _cvpt_3019;   // oc8051_tb.v(104)
    output _cvpt_3020;   // oc8051_tb.v(104)
    output _cvpt_3021;   // oc8051_tb.v(104)
    output _cvpt_3022;   // oc8051_tb.v(104)
    output _cvpt_3023;   // oc8051_tb.v(104)
    output _cvpt_3024;   // oc8051_tb.v(104)
    output _cvpt_3025;   // oc8051_tb.v(104)
    output _cvpt_3026;   // oc8051_tb.v(104)
    output _cvpt_3027;   // oc8051_tb.v(104)
    output _cvpt_3028;   // oc8051_tb.v(104)
    output _cvpt_3029;   // oc8051_tb.v(104)
    output _cvpt_3030;   // oc8051_tb.v(104)
    output _cvpt_3031;   // oc8051_tb.v(104)
    output _cvpt_3032;   // oc8051_tb.v(104)
    output _cvpt_3033;   // oc8051_tb.v(104)
    output _cvpt_3034;   // oc8051_tb.v(104)
    output _cvpt_3035;   // oc8051_tb.v(104)
    output _cvpt_3036;   // oc8051_tb.v(104)
    output _cvpt_3037;   // oc8051_tb.v(104)
    output _cvpt_3038;   // oc8051_tb.v(104)
    output _cvpt_3039;   // oc8051_tb.v(104)
    output _cvpt_3040;   // oc8051_tb.v(104)
    output _cvpt_3041;   // oc8051_tb.v(104)
    output _cvpt_3042;   // oc8051_tb.v(104)
    output _cvpt_3043;   // oc8051_tb.v(104)
    output _cvpt_3044;   // oc8051_tb.v(104)
    output _cvpt_3045;   // oc8051_tb.v(104)
    output _cvpt_3046;   // oc8051_tb.v(104)
    output _cvpt_3047;   // oc8051_tb.v(104)
    output _cvpt_3048;   // oc8051_tb.v(104)
    output _cvpt_3049;   // oc8051_tb.v(104)
    output _cvpt_3050;   // oc8051_tb.v(104)
    output _cvpt_3051;   // oc8051_tb.v(104)
    output _cvpt_3052;   // oc8051_tb.v(104)
    output _cvpt_3053;   // oc8051_tb.v(104)
    output _cvpt_3054;   // oc8051_tb.v(104)
    output _cvpt_3055;   // oc8051_tb.v(104)
    output _cvpt_3056;   // oc8051_tb.v(104)
    output _cvpt_3057;   // oc8051_tb.v(104)
    output _cvpt_3058;   // oc8051_tb.v(104)
    output _cvpt_3059;   // oc8051_tb.v(104)
    output _cvpt_3060;   // oc8051_tb.v(104)
    output _cvpt_3061;   // oc8051_tb.v(104)
    output _cvpt_3062;   // oc8051_tb.v(104)
    output _cvpt_3063;   // oc8051_tb.v(104)
    output _cvpt_3064;   // oc8051_tb.v(104)
    output _cvpt_3065;   // oc8051_tb.v(104)
    output _cvpt_3066;   // oc8051_tb.v(104)
    output _cvpt_3067;   // oc8051_tb.v(104)
    output _cvpt_3068;   // oc8051_tb.v(104)
    output _cvpt_3069;   // oc8051_tb.v(104)
    output _cvpt_3070;   // oc8051_tb.v(104)
    output _cvpt_3071;   // oc8051_tb.v(104)
    output _cvpt_3072;   // oc8051_tb.v(104)
    output _cvpt_3073;   // oc8051_tb.v(104)
    output _cvpt_3074;   // oc8051_tb.v(104)
    output _cvpt_3075;   // oc8051_tb.v(104)
    output _cvpt_3076;   // oc8051_tb.v(104)
    output _cvpt_3077;   // oc8051_tb.v(104)
    output _cvpt_3078;   // oc8051_tb.v(104)
    output _cvpt_3079;   // oc8051_tb.v(104)
    output _cvpt_3080;   // oc8051_tb.v(104)
    output _cvpt_3081;   // oc8051_tb.v(104)
    output _cvpt_3082;   // oc8051_tb.v(104)
    output _cvpt_3083;   // oc8051_tb.v(104)
    output _cvpt_3084;   // oc8051_tb.v(104)
    output _cvpt_3085;   // oc8051_tb.v(104)
    output _cvpt_3086;   // oc8051_tb.v(104)
    output _cvpt_3087;   // oc8051_tb.v(104)
    output _cvpt_3088;   // oc8051_tb.v(104)
    output _cvpt_3089;   // oc8051_tb.v(104)
    output _cvpt_3090;   // oc8051_tb.v(104)
    output _cvpt_3091;   // oc8051_tb.v(104)
    output _cvpt_3092;   // oc8051_tb.v(104)
    output _cvpt_3093;   // oc8051_tb.v(104)
    output _cvpt_3094;   // oc8051_tb.v(104)
    output _cvpt_3095;   // oc8051_tb.v(104)
    output _cvpt_3096;   // oc8051_tb.v(104)
    output _cvpt_3097;   // oc8051_tb.v(104)
    output _cvpt_3098;   // oc8051_tb.v(104)
    output _cvpt_3099;   // oc8051_tb.v(104)
    output _cvpt_3100;   // oc8051_tb.v(104)
    output _cvpt_3101;   // oc8051_tb.v(104)
    output _cvpt_3102;   // oc8051_tb.v(104)
    output _cvpt_3103;   // oc8051_tb.v(104)
    output _cvpt_3104;   // oc8051_tb.v(104)
    output _cvpt_3105;   // oc8051_tb.v(104)
    output _cvpt_3106;   // oc8051_tb.v(104)
    output _cvpt_3107;   // oc8051_tb.v(104)
    output _cvpt_3108;   // oc8051_tb.v(104)
    output _cvpt_3109;   // oc8051_tb.v(104)
    output _cvpt_3110;   // oc8051_tb.v(104)
    output _cvpt_3111;   // oc8051_tb.v(104)
    output _cvpt_3112;   // oc8051_tb.v(104)
    output _cvpt_3113;   // oc8051_tb.v(104)
    output _cvpt_3114;   // oc8051_tb.v(104)
    output _cvpt_3115;   // oc8051_tb.v(104)
    output _cvpt_3116;   // oc8051_tb.v(104)
    output _cvpt_3117;   // oc8051_tb.v(104)
    output _cvpt_3118;   // oc8051_tb.v(104)
    output _cvpt_3119;   // oc8051_tb.v(104)
    output _cvpt_3120;   // oc8051_tb.v(104)
    output _cvpt_3121;   // oc8051_tb.v(104)
    output _cvpt_3122;   // oc8051_tb.v(104)
    output _cvpt_3123;   // oc8051_tb.v(104)
    output _cvpt_3124;   // oc8051_tb.v(104)
    output _cvpt_3125;   // oc8051_tb.v(104)
    output _cvpt_3126;   // oc8051_tb.v(104)
    output _cvpt_3127;   // oc8051_tb.v(104)
    output _cvpt_3128;   // oc8051_tb.v(104)
    output _cvpt_3129;   // oc8051_tb.v(104)
    output _cvpt_3130;   // oc8051_tb.v(104)
    output _cvpt_3131;   // oc8051_tb.v(104)
    output _cvpt_3132;   // oc8051_tb.v(104)
    output _cvpt_3133;   // oc8051_tb.v(104)
    output _cvpt_3134;   // oc8051_tb.v(104)
    output _cvpt_3135;   // oc8051_tb.v(104)
    output _cvpt_3136;   // oc8051_tb.v(104)
    output _cvpt_3137;   // oc8051_tb.v(104)
    output _cvpt_3138;   // oc8051_tb.v(104)
    output _cvpt_3139;   // oc8051_tb.v(104)
    output _cvpt_3140;   // oc8051_tb.v(104)
    output _cvpt_3141;   // oc8051_tb.v(104)
    output _cvpt_3142;   // oc8051_tb.v(104)
    output _cvpt_3143;   // oc8051_tb.v(104)
    output _cvpt_3144;   // oc8051_tb.v(104)
    output _cvpt_3145;   // oc8051_tb.v(104)
    output _cvpt_3146;   // oc8051_tb.v(104)
    output _cvpt_3147;   // oc8051_tb.v(104)
    output _cvpt_3148;   // oc8051_tb.v(104)
    output _cvpt_3149;   // oc8051_tb.v(104)
    output _cvpt_3150;   // oc8051_tb.v(104)
    output _cvpt_3151;   // oc8051_tb.v(104)
    output _cvpt_3152;   // oc8051_tb.v(104)
    output _cvpt_3153;   // oc8051_tb.v(104)
    output _cvpt_3154;   // oc8051_tb.v(104)
    output _cvpt_3155;   // oc8051_tb.v(104)
    output _cvpt_3156;   // oc8051_tb.v(104)
    output _cvpt_3157;   // oc8051_tb.v(104)
    output _cvpt_3158;   // oc8051_tb.v(104)
    output _cvpt_3159;   // oc8051_tb.v(104)
    output _cvpt_3160;   // oc8051_tb.v(104)
    output _cvpt_3161;   // oc8051_tb.v(104)
    output _cvpt_3162;   // oc8051_tb.v(104)
    output _cvpt_3163;   // oc8051_tb.v(104)
    output _cvpt_3164;   // oc8051_tb.v(104)
    output _cvpt_3165;   // oc8051_tb.v(104)
    output _cvpt_3166;   // oc8051_tb.v(104)
    output _cvpt_3167;   // oc8051_tb.v(104)
    output _cvpt_3168;   // oc8051_tb.v(104)
    output _cvpt_3169;   // oc8051_tb.v(104)
    output _cvpt_3170;   // oc8051_tb.v(104)
    output _cvpt_3171;   // oc8051_tb.v(104)
    output _cvpt_3172;   // oc8051_tb.v(104)
    output _cvpt_3173;   // oc8051_tb.v(104)
    output _cvpt_3174;   // oc8051_tb.v(104)
    output _cvpt_3175;   // oc8051_tb.v(104)
    output _cvpt_3176;   // oc8051_tb.v(104)
    output _cvpt_3177;   // oc8051_tb.v(104)
    output _cvpt_3178;   // oc8051_tb.v(104)
    output _cvpt_3179;   // oc8051_tb.v(104)
    output _cvpt_3180;   // oc8051_tb.v(104)
    output _cvpt_3181;   // oc8051_tb.v(104)
    output _cvpt_3182;   // oc8051_tb.v(104)
    output _cvpt_3183;   // oc8051_tb.v(104)
    output _cvpt_3184;   // oc8051_tb.v(104)
    output _cvpt_3185;   // oc8051_tb.v(104)
    output _cvpt_3186;   // oc8051_tb.v(104)
    output _cvpt_3187;   // oc8051_tb.v(104)
    output _cvpt_3188;   // oc8051_tb.v(104)
    output _cvpt_3189;   // oc8051_tb.v(104)
    output _cvpt_3190;   // oc8051_tb.v(104)
    output _cvpt_3191;   // oc8051_tb.v(104)
    output _cvpt_3192;   // oc8051_tb.v(104)
    output _cvpt_3193;   // oc8051_tb.v(104)
    output _cvpt_3194;   // oc8051_tb.v(104)
    output _cvpt_3195;   // oc8051_tb.v(104)
    output _cvpt_3196;   // oc8051_tb.v(104)
    output _cvpt_3197;   // oc8051_tb.v(104)
    output _cvpt_3198;   // oc8051_tb.v(104)
    output _cvpt_3199;   // oc8051_tb.v(104)
    output _cvpt_3200;   // oc8051_tb.v(104)
    output _cvpt_3201;   // oc8051_tb.v(104)
    output _cvpt_3202;   // oc8051_tb.v(104)
    output _cvpt_3203;   // oc8051_tb.v(104)
    output _cvpt_3204;   // oc8051_tb.v(104)
    output _cvpt_3205;   // oc8051_tb.v(104)
    output _cvpt_3206;   // oc8051_tb.v(104)
    output _cvpt_3207;   // oc8051_tb.v(104)
    output _cvpt_3208;   // oc8051_tb.v(104)
    output _cvpt_3209;   // oc8051_tb.v(104)
    output _cvpt_3210;   // oc8051_tb.v(104)
    output _cvpt_3211;   // oc8051_tb.v(104)
    output _cvpt_3212;   // oc8051_tb.v(104)
    output _cvpt_3213;   // oc8051_tb.v(104)
    output _cvpt_3214;   // oc8051_tb.v(104)
    output _cvpt_3215;   // oc8051_tb.v(104)
    output _cvpt_3216;   // oc8051_tb.v(104)
    output _cvpt_3217;   // oc8051_tb.v(104)
    output _cvpt_3218;   // oc8051_tb.v(104)
    output _cvpt_3219;   // oc8051_tb.v(104)
    output _cvpt_3220;   // oc8051_tb.v(104)
    output _cvpt_3221;   // oc8051_tb.v(104)
    output _cvpt_3222;   // oc8051_tb.v(104)
    output _cvpt_3223;   // oc8051_tb.v(104)
    output _cvpt_3224;   // oc8051_tb.v(104)
    output _cvpt_3225;   // oc8051_tb.v(104)
    output _cvpt_3226;   // oc8051_tb.v(104)
    output _cvpt_3227;   // oc8051_tb.v(104)
    output _cvpt_3228;   // oc8051_tb.v(104)
    output _cvpt_3229;   // oc8051_tb.v(104)
    output _cvpt_3230;   // oc8051_tb.v(104)
    output _cvpt_3231;   // oc8051_tb.v(104)
    output _cvpt_3232;   // oc8051_tb.v(104)
    output _cvpt_3233;   // oc8051_tb.v(104)
    output _cvpt_3234;   // oc8051_tb.v(104)
    output _cvpt_3235;   // oc8051_tb.v(104)
    output _cvpt_3236;   // oc8051_tb.v(104)
    output _cvpt_3237;   // oc8051_tb.v(104)
    output _cvpt_3238;   // oc8051_tb.v(104)
    output _cvpt_3239;   // oc8051_tb.v(104)
    output _cvpt_3240;   // oc8051_tb.v(104)
    output _cvpt_3241;   // oc8051_tb.v(104)
    output _cvpt_3242;   // oc8051_tb.v(104)
    output _cvpt_3243;   // oc8051_tb.v(104)
    output _cvpt_3244;   // oc8051_tb.v(104)
    output _cvpt_3245;   // oc8051_tb.v(104)
    output _cvpt_3246;   // oc8051_tb.v(104)
    output _cvpt_3247;   // oc8051_tb.v(104)
    output _cvpt_3248;   // oc8051_tb.v(104)
    output _cvpt_3249;   // oc8051_tb.v(104)
    output _cvpt_3250;   // oc8051_tb.v(104)
    output _cvpt_3251;   // oc8051_tb.v(104)
    output _cvpt_3252;   // oc8051_tb.v(104)
    output _cvpt_3253;   // oc8051_tb.v(104)
    output _cvpt_3254;   // oc8051_tb.v(104)
    output _cvpt_3255;   // oc8051_tb.v(104)
    output _cvpt_3256;   // oc8051_tb.v(104)
    output _cvpt_3257;   // oc8051_tb.v(104)
    output _cvpt_3258;   // oc8051_tb.v(104)
    output _cvpt_3259;   // oc8051_tb.v(104)
    output _cvpt_3260;   // oc8051_tb.v(104)
    output _cvpt_3261;   // oc8051_tb.v(104)
    output _cvpt_3262;   // oc8051_tb.v(104)
    output _cvpt_3263;   // oc8051_tb.v(104)
    output _cvpt_3264;   // oc8051_tb.v(104)
    output _cvpt_3265;   // oc8051_tb.v(104)
    output _cvpt_3266;   // oc8051_tb.v(104)
    output _cvpt_3267;   // oc8051_tb.v(104)
    output _cvpt_3268;   // oc8051_tb.v(104)
    output _cvpt_3269;   // oc8051_tb.v(104)
    output _cvpt_3270;   // oc8051_tb.v(104)
    output _cvpt_3271;   // oc8051_tb.v(104)
    output _cvpt_3272;   // oc8051_tb.v(104)
    output _cvpt_3273;   // oc8051_tb.v(104)
    output _cvpt_3274;   // oc8051_tb.v(104)
    output _cvpt_3275;   // oc8051_tb.v(104)
    output _cvpt_3276;   // oc8051_tb.v(104)
    output _cvpt_3277;   // oc8051_tb.v(104)
    output _cvpt_3278;   // oc8051_tb.v(104)
    output _cvpt_3279;   // oc8051_tb.v(104)
    output _cvpt_3280;   // oc8051_tb.v(104)
    output _cvpt_3281;   // oc8051_tb.v(104)
    output _cvpt_3282;   // oc8051_tb.v(104)
    output _cvpt_3283;   // oc8051_tb.v(104)
    output _cvpt_3284;   // oc8051_tb.v(104)
    output _cvpt_3285;   // oc8051_tb.v(104)
    output _cvpt_3286;   // oc8051_tb.v(104)
    output _cvpt_3287;   // oc8051_tb.v(104)
    output _cvpt_3288;   // oc8051_tb.v(104)
    output _cvpt_3289;   // oc8051_tb.v(104)
    output _cvpt_3290;   // oc8051_tb.v(104)
    output _cvpt_3291;   // oc8051_tb.v(104)
    output _cvpt_3292;   // oc8051_tb.v(104)
    output _cvpt_3293;   // oc8051_tb.v(104)
    output _cvpt_3294;   // oc8051_tb.v(104)
    output _cvpt_3295;   // oc8051_tb.v(104)
    output _cvpt_3296;   // oc8051_tb.v(104)
    output _cvpt_3297;   // oc8051_tb.v(104)
    output _cvpt_3298;   // oc8051_tb.v(104)
    output _cvpt_3299;   // oc8051_tb.v(104)
    output _cvpt_3300;   // oc8051_tb.v(104)
    output _cvpt_3301;   // oc8051_tb.v(104)
    output _cvpt_3302;   // oc8051_tb.v(104)
    output _cvpt_3303;   // oc8051_tb.v(104)
    output _cvpt_3304;   // oc8051_tb.v(104)
    output _cvpt_3305;   // oc8051_tb.v(104)
    output _cvpt_3306;   // oc8051_tb.v(104)
    output _cvpt_3307;   // oc8051_tb.v(104)
    output _cvpt_3308;   // oc8051_tb.v(104)
    output _cvpt_3309;   // oc8051_tb.v(104)
    output _cvpt_3310;   // oc8051_tb.v(104)
    output _cvpt_3311;   // oc8051_tb.v(104)
    output _cvpt_3312;   // oc8051_tb.v(104)
    output _cvpt_3313;   // oc8051_tb.v(104)
    output _cvpt_3314;   // oc8051_tb.v(104)
    output _cvpt_3315;   // oc8051_tb.v(104)
    output _cvpt_3316;   // oc8051_tb.v(104)
    output _cvpt_3317;   // oc8051_tb.v(104)
    output _cvpt_3318;   // oc8051_tb.v(104)
    output _cvpt_3319;   // oc8051_tb.v(104)
    output _cvpt_3320;   // oc8051_tb.v(104)
    output _cvpt_3321;   // oc8051_tb.v(104)
    output _cvpt_3322;   // oc8051_tb.v(104)
    output _cvpt_3323;   // oc8051_tb.v(104)
    output _cvpt_3324;   // oc8051_tb.v(104)
    output _cvpt_3325;   // oc8051_tb.v(104)
    output _cvpt_3326;   // oc8051_tb.v(104)
    output _cvpt_3327;   // oc8051_tb.v(104)
    output _cvpt_3328;   // oc8051_tb.v(104)
    output _cvpt_3329;   // oc8051_tb.v(104)
    output _cvpt_3330;   // oc8051_tb.v(104)
    output _cvpt_3331;   // oc8051_tb.v(104)
    output _cvpt_3332;   // oc8051_tb.v(104)
    output _cvpt_3333;   // oc8051_tb.v(104)
    output _cvpt_3334;   // oc8051_tb.v(104)
    output _cvpt_3335;   // oc8051_tb.v(104)
    output _cvpt_3336;   // oc8051_tb.v(104)
    output _cvpt_3337;   // oc8051_tb.v(104)
    output _cvpt_3338;   // oc8051_tb.v(104)
    output _cvpt_3339;   // oc8051_tb.v(104)
    output _cvpt_3340;   // oc8051_tb.v(104)
    output _cvpt_3341;   // oc8051_tb.v(104)
    output _cvpt_3342;   // oc8051_tb.v(104)
    output _cvpt_3343;   // oc8051_tb.v(104)
    output _cvpt_3344;   // oc8051_tb.v(104)
    output _cvpt_3345;   // oc8051_tb.v(104)
    output _cvpt_3346;   // oc8051_tb.v(104)
    output _cvpt_3347;   // oc8051_tb.v(104)
    output _cvpt_3348;   // oc8051_tb.v(104)
    output _cvpt_3349;   // oc8051_tb.v(104)
    output _cvpt_3350;   // oc8051_tb.v(104)
    output _cvpt_3351;   // oc8051_tb.v(104)
    output _cvpt_3352;   // oc8051_tb.v(104)
    output _cvpt_3353;   // oc8051_tb.v(104)
    output _cvpt_3354;   // oc8051_tb.v(104)
    output _cvpt_3355;   // oc8051_tb.v(104)
    output _cvpt_3356;   // oc8051_tb.v(104)
    output _cvpt_3357;   // oc8051_tb.v(104)
    output _cvpt_3358;   // oc8051_tb.v(104)
    output _cvpt_3359;   // oc8051_tb.v(104)
    output _cvpt_3360;   // oc8051_tb.v(104)
    output _cvpt_3361;   // oc8051_tb.v(104)
    output _cvpt_3362;   // oc8051_tb.v(104)
    output _cvpt_3363;   // oc8051_tb.v(104)
    output _cvpt_3364;   // oc8051_tb.v(104)
    output _cvpt_3365;   // oc8051_tb.v(104)
    output _cvpt_3366;   // oc8051_tb.v(104)
    output _cvpt_3367;   // oc8051_tb.v(104)
    output _cvpt_3368;   // oc8051_tb.v(104)
    output _cvpt_3369;   // oc8051_tb.v(104)
    output _cvpt_3370;   // oc8051_tb.v(104)
    output _cvpt_3371;   // oc8051_tb.v(104)
    output _cvpt_3372;   // oc8051_tb.v(104)
    output _cvpt_3373;   // oc8051_tb.v(104)
    output _cvpt_3374;   // oc8051_tb.v(104)
    output _cvpt_3375;   // oc8051_tb.v(104)
    output _cvpt_3376;   // oc8051_tb.v(104)
    output _cvpt_3377;   // oc8051_tb.v(104)
    output _cvpt_3378;   // oc8051_tb.v(104)
    output _cvpt_3379;   // oc8051_tb.v(104)
    output _cvpt_3380;   // oc8051_tb.v(104)
    output _cvpt_3381;   // oc8051_tb.v(104)
    output _cvpt_3382;   // oc8051_tb.v(104)
    output _cvpt_3383;   // oc8051_tb.v(104)
    output _cvpt_3384;   // oc8051_tb.v(104)
    output _cvpt_3385;   // oc8051_tb.v(104)
    output _cvpt_3386;   // oc8051_tb.v(104)
    output _cvpt_3387;   // oc8051_tb.v(104)
    output _cvpt_3388;   // oc8051_tb.v(104)
    output _cvpt_3389;   // oc8051_tb.v(104)
    output _cvpt_3390;   // oc8051_tb.v(104)
    output _cvpt_3391;   // oc8051_tb.v(104)
    output _cvpt_3392;   // oc8051_tb.v(104)
    output _cvpt_3393;   // oc8051_tb.v(104)
    output _cvpt_3394;   // oc8051_tb.v(104)
    output _cvpt_3395;   // oc8051_tb.v(104)
    output _cvpt_3396;   // oc8051_tb.v(104)
    output _cvpt_3397;   // oc8051_tb.v(104)
    output _cvpt_3398;   // oc8051_tb.v(104)
    output _cvpt_3399;   // oc8051_tb.v(104)
    output _cvpt_3400;   // oc8051_tb.v(104)
    output _cvpt_3401;   // oc8051_tb.v(104)
    output _cvpt_3402;   // oc8051_tb.v(104)
    output _cvpt_3403;   // oc8051_tb.v(104)
    output _cvpt_3404;   // oc8051_tb.v(104)
    output _cvpt_3405;   // oc8051_tb.v(104)
    output _cvpt_3406;   // oc8051_tb.v(104)
    output _cvpt_3407;   // oc8051_tb.v(104)
    output _cvpt_3408;   // oc8051_tb.v(104)
    output _cvpt_3409;   // oc8051_tb.v(104)
    output _cvpt_3410;   // oc8051_tb.v(104)
    output _cvpt_3411;   // oc8051_tb.v(104)
    output _cvpt_3412;   // oc8051_tb.v(104)
    output _cvpt_3413;   // oc8051_tb.v(104)
    output _cvpt_3414;   // oc8051_tb.v(104)
    output _cvpt_3415;   // oc8051_tb.v(104)
    output _cvpt_3416;   // oc8051_tb.v(104)
    output _cvpt_3417;   // oc8051_tb.v(104)
    output _cvpt_3418;   // oc8051_tb.v(104)
    output _cvpt_3419;   // oc8051_tb.v(104)
    output _cvpt_3420;   // oc8051_tb.v(104)
    output _cvpt_3421;   // oc8051_tb.v(104)
    output _cvpt_3422;   // oc8051_tb.v(104)
    output _cvpt_3423;   // oc8051_tb.v(104)
    output _cvpt_3424;   // oc8051_tb.v(104)
    output _cvpt_3425;   // oc8051_tb.v(104)
    output _cvpt_3426;   // oc8051_tb.v(104)
    output _cvpt_3427;   // oc8051_tb.v(104)
    output _cvpt_3428;   // oc8051_tb.v(104)
    output _cvpt_3429;   // oc8051_tb.v(104)
    output _cvpt_3430;   // oc8051_tb.v(104)
    output _cvpt_3431;   // oc8051_tb.v(104)
    output _cvpt_3432;   // oc8051_tb.v(104)
    output _cvpt_3433;   // oc8051_tb.v(104)
    output _cvpt_3434;   // oc8051_tb.v(104)
    output _cvpt_3435;   // oc8051_tb.v(104)
    output _cvpt_3436;   // oc8051_tb.v(104)
    output _cvpt_3437;   // oc8051_tb.v(104)
    output _cvpt_3438;   // oc8051_tb.v(104)
    output _cvpt_3439;   // oc8051_tb.v(104)
    output _cvpt_3440;   // oc8051_tb.v(104)
    output _cvpt_3441;   // oc8051_tb.v(104)
    output _cvpt_3442;   // oc8051_tb.v(104)
    output _cvpt_3443;   // oc8051_tb.v(104)
    output _cvpt_3444;   // oc8051_tb.v(104)
    output _cvpt_3445;   // oc8051_tb.v(104)
    output _cvpt_3446;   // oc8051_tb.v(104)
    output _cvpt_3447;   // oc8051_tb.v(104)
    output _cvpt_3448;   // oc8051_tb.v(104)
    output _cvpt_3449;   // oc8051_tb.v(104)
    output _cvpt_3450;   // oc8051_tb.v(104)
    output _cvpt_3451;   // oc8051_tb.v(104)
    output _cvpt_3452;   // oc8051_tb.v(104)
    output _cvpt_3453;   // oc8051_tb.v(104)
    output _cvpt_3454;   // oc8051_tb.v(104)
    output _cvpt_3455;   // oc8051_tb.v(104)
    output _cvpt_3456;   // oc8051_tb.v(104)
    output _cvpt_3457;   // oc8051_tb.v(104)
    output _cvpt_3458;   // oc8051_tb.v(104)
    output _cvpt_3459;   // oc8051_tb.v(104)
    output _cvpt_3460;   // oc8051_tb.v(104)
    output _cvpt_3461;   // oc8051_tb.v(104)
    output _cvpt_3462;   // oc8051_tb.v(104)
    output _cvpt_3463;   // oc8051_tb.v(104)
    output _cvpt_3464;   // oc8051_tb.v(104)
    output _cvpt_3465;   // oc8051_tb.v(104)
    output _cvpt_3466;   // oc8051_tb.v(104)
    output _cvpt_3467;   // oc8051_tb.v(104)
    output _cvpt_3468;   // oc8051_tb.v(104)
    output _cvpt_3469;   // oc8051_tb.v(104)
    output _cvpt_3470;   // oc8051_tb.v(104)
    output _cvpt_3471;   // oc8051_tb.v(104)
    output _cvpt_3472;   // oc8051_tb.v(104)
    output _cvpt_3473;   // oc8051_tb.v(104)
    output _cvpt_3474;   // oc8051_tb.v(104)
    output _cvpt_3475;   // oc8051_tb.v(104)
    output _cvpt_3476;   // oc8051_tb.v(104)
    output _cvpt_3477;   // oc8051_tb.v(104)
    output _cvpt_3478;   // oc8051_tb.v(104)
    output _cvpt_3479;   // oc8051_tb.v(104)
    output _cvpt_3480;   // oc8051_tb.v(104)
    output _cvpt_3481;   // oc8051_tb.v(104)
    output _cvpt_3482;   // oc8051_tb.v(104)
    output _cvpt_3483;   // oc8051_tb.v(104)
    output _cvpt_3484;   // oc8051_tb.v(104)
    output _cvpt_3485;   // oc8051_tb.v(104)
    output _cvpt_3486;   // oc8051_tb.v(104)
    output _cvpt_3487;   // oc8051_tb.v(104)
    output _cvpt_3488;   // oc8051_tb.v(104)
    output _cvpt_3489;   // oc8051_tb.v(104)
    output _cvpt_3490;   // oc8051_tb.v(104)
    output _cvpt_3491;   // oc8051_tb.v(104)
    output _cvpt_3492;   // oc8051_tb.v(104)
    output _cvpt_3493;   // oc8051_tb.v(104)
    output _cvpt_3494;   // oc8051_tb.v(104)
    output _cvpt_3495;   // oc8051_tb.v(104)
    output _cvpt_3496;   // oc8051_tb.v(104)
    output _cvpt_3497;   // oc8051_tb.v(104)
    output _cvpt_3498;   // oc8051_tb.v(104)
    output _cvpt_3499;   // oc8051_tb.v(104)
    output _cvpt_3500;   // oc8051_tb.v(104)
    output _cvpt_3501;   // oc8051_tb.v(104)
    output _cvpt_3502;   // oc8051_tb.v(104)
    output _cvpt_3503;   // oc8051_tb.v(104)
    output _cvpt_3504;   // oc8051_tb.v(104)
    output _cvpt_3505;   // oc8051_tb.v(104)
    output _cvpt_3506;   // oc8051_tb.v(104)
    output _cvpt_3507;   // oc8051_tb.v(104)
    output _cvpt_3508;   // oc8051_tb.v(104)
    output _cvpt_3509;   // oc8051_tb.v(104)
    output _cvpt_3510;   // oc8051_tb.v(104)
    output _cvpt_3511;   // oc8051_tb.v(104)
    output _cvpt_3512;   // oc8051_tb.v(104)
    output _cvpt_3513;   // oc8051_tb.v(104)
    output _cvpt_3514;   // oc8051_tb.v(104)
    output _cvpt_3515;   // oc8051_tb.v(104)
    output _cvpt_3516;   // oc8051_tb.v(104)
    output _cvpt_3517;   // oc8051_tb.v(104)
    output _cvpt_3518;   // oc8051_tb.v(104)
    output _cvpt_3519;   // oc8051_tb.v(104)
    output _cvpt_3520;   // oc8051_tb.v(104)
    output _cvpt_3521;   // oc8051_tb.v(104)
    output _cvpt_3522;   // oc8051_tb.v(104)
    output _cvpt_3523;   // oc8051_tb.v(104)
    output _cvpt_3524;   // oc8051_tb.v(104)
    output _cvpt_3525;   // oc8051_tb.v(104)
    output _cvpt_3526;   // oc8051_tb.v(104)
    output _cvpt_3527;   // oc8051_tb.v(104)
    output _cvpt_3528;   // oc8051_tb.v(104)
    output _cvpt_3529;   // oc8051_tb.v(104)
    output _cvpt_3530;   // oc8051_tb.v(104)
    output _cvpt_3531;   // oc8051_tb.v(104)
    output _cvpt_3532;   // oc8051_tb.v(104)
    output _cvpt_3533;   // oc8051_tb.v(104)
    output _cvpt_3534;   // oc8051_tb.v(104)
    output _cvpt_3535;   // oc8051_tb.v(104)
    output _cvpt_3536;   // oc8051_tb.v(104)
    output _cvpt_3537;   // oc8051_tb.v(104)
    output _cvpt_3538;   // oc8051_tb.v(104)
    output _cvpt_3539;   // oc8051_tb.v(104)
    output _cvpt_3540;   // oc8051_tb.v(104)
    output _cvpt_3541;   // oc8051_tb.v(104)
    output _cvpt_3542;   // oc8051_tb.v(104)
    output _cvpt_3543;   // oc8051_tb.v(104)
    output _cvpt_3544;   // oc8051_tb.v(104)
    output _cvpt_3545;   // oc8051_tb.v(104)
    output _cvpt_3546;   // oc8051_tb.v(104)
    output _cvpt_3547;   // oc8051_tb.v(104)
    output _cvpt_3548;   // oc8051_tb.v(104)
    output _cvpt_3549;   // oc8051_tb.v(104)
    output _cvpt_3550;   // oc8051_tb.v(104)
    output _cvpt_3551;   // oc8051_tb.v(104)
    output _cvpt_3552;   // oc8051_tb.v(104)
    output _cvpt_3553;   // oc8051_tb.v(104)
    output _cvpt_3554;   // oc8051_tb.v(104)
    output _cvpt_3555;   // oc8051_tb.v(104)
    output _cvpt_3556;   // oc8051_tb.v(104)
    output _cvpt_3557;   // oc8051_tb.v(104)
    output _cvpt_3558;   // oc8051_tb.v(104)
    output _cvpt_3559;   // oc8051_tb.v(104)
    output _cvpt_3560;   // oc8051_tb.v(104)
    output _cvpt_3561;   // oc8051_tb.v(104)
    output _cvpt_3562;   // oc8051_tb.v(104)
    output _cvpt_3563;   // oc8051_tb.v(104)
    output _cvpt_3564;   // oc8051_tb.v(104)
    output _cvpt_3565;   // oc8051_tb.v(104)
    output _cvpt_3566;   // oc8051_tb.v(104)
    output _cvpt_3567;   // oc8051_tb.v(104)
    output _cvpt_3568;   // oc8051_tb.v(104)
    output _cvpt_3569;   // oc8051_tb.v(104)
    output _cvpt_3570;   // oc8051_tb.v(104)
    output _cvpt_3571;   // oc8051_tb.v(104)
    output _cvpt_3572;   // oc8051_tb.v(104)
    output _cvpt_3573;   // oc8051_tb.v(104)
    output _cvpt_3574;   // oc8051_tb.v(104)
    output _cvpt_3575;   // oc8051_tb.v(104)
    output _cvpt_3576;   // oc8051_tb.v(104)
    output _cvpt_3577;   // oc8051_tb.v(104)
    output _cvpt_3578;   // oc8051_tb.v(104)
    output _cvpt_3579;   // oc8051_tb.v(104)
    output _cvpt_3580;   // oc8051_tb.v(104)
    output _cvpt_3581;   // oc8051_tb.v(104)
    output _cvpt_3582;   // oc8051_tb.v(104)
    output _cvpt_3583;   // oc8051_tb.v(104)
    output _cvpt_3584;   // oc8051_tb.v(104)
    output _cvpt_3585;   // oc8051_tb.v(104)
    output _cvpt_3586;   // oc8051_tb.v(104)
    output _cvpt_3587;   // oc8051_tb.v(104)
    output _cvpt_3588;   // oc8051_tb.v(104)
    output _cvpt_3589;   // oc8051_tb.v(104)
    output _cvpt_3590;   // oc8051_tb.v(104)
    output _cvpt_3591;   // oc8051_tb.v(104)
    output _cvpt_3592;   // oc8051_tb.v(104)
    output _cvpt_3593;   // oc8051_tb.v(104)
    output _cvpt_3594;   // oc8051_tb.v(104)
    output _cvpt_3595;   // oc8051_tb.v(104)
    output _cvpt_3596;   // oc8051_tb.v(104)
    output _cvpt_3597;   // oc8051_tb.v(104)
    output _cvpt_3598;   // oc8051_tb.v(104)
    output _cvpt_3599;   // oc8051_tb.v(104)
    output _cvpt_3600;   // oc8051_tb.v(104)
    output _cvpt_3601;   // oc8051_tb.v(104)
    output _cvpt_3602;   // oc8051_tb.v(104)
    output _cvpt_3603;   // oc8051_tb.v(104)
    output _cvpt_3604;   // oc8051_tb.v(104)
    output _cvpt_3605;   // oc8051_tb.v(104)
    output _cvpt_3606;   // oc8051_tb.v(104)
    output _cvpt_3607;   // oc8051_tb.v(104)
    output _cvpt_3608;   // oc8051_tb.v(104)
    output _cvpt_3609;   // oc8051_tb.v(104)
    output _cvpt_3610;   // oc8051_tb.v(104)
    output _cvpt_3611;   // oc8051_tb.v(104)
    output _cvpt_3612;   // oc8051_tb.v(104)
    output _cvpt_3613;   // oc8051_tb.v(104)
    output _cvpt_3614;   // oc8051_tb.v(104)
    output _cvpt_3615;   // oc8051_tb.v(104)
    output _cvpt_3616;   // oc8051_tb.v(104)
    output _cvpt_3617;   // oc8051_tb.v(104)
    output _cvpt_3618;   // oc8051_tb.v(104)
    output _cvpt_3619;   // oc8051_tb.v(104)
    output _cvpt_3620;   // oc8051_tb.v(104)
    output _cvpt_3621;   // oc8051_tb.v(104)
    output _cvpt_3622;   // oc8051_tb.v(104)
    output _cvpt_3623;   // oc8051_tb.v(104)
    output _cvpt_3624;   // oc8051_tb.v(104)
    output _cvpt_3625;   // oc8051_tb.v(104)
    output _cvpt_3626;   // oc8051_tb.v(104)
    output _cvpt_3627;   // oc8051_tb.v(104)
    output _cvpt_3628;   // oc8051_tb.v(104)
    output _cvpt_3629;   // oc8051_tb.v(104)
    output _cvpt_3630;   // oc8051_tb.v(104)
    output _cvpt_3631;   // oc8051_tb.v(104)
    output _cvpt_3632;   // oc8051_tb.v(104)
    output _cvpt_3633;   // oc8051_tb.v(104)
    output _cvpt_3634;   // oc8051_tb.v(104)
    output _cvpt_3635;   // oc8051_tb.v(104)
    output _cvpt_3636;   // oc8051_tb.v(104)
    output _cvpt_3637;   // oc8051_tb.v(104)
    output _cvpt_3638;   // oc8051_tb.v(104)
    output _cvpt_3639;   // oc8051_tb.v(104)
    output _cvpt_3640;   // oc8051_tb.v(104)
    output _cvpt_3641;   // oc8051_tb.v(104)
    output _cvpt_3642;   // oc8051_tb.v(104)
    output _cvpt_3643;   // oc8051_tb.v(104)
    output _cvpt_3644;   // oc8051_tb.v(104)
    output _cvpt_3645;   // oc8051_tb.v(104)
    output _cvpt_3646;   // oc8051_tb.v(104)
    output _cvpt_3647;   // oc8051_tb.v(104)
    output _cvpt_3648;   // oc8051_tb.v(104)
    output _cvpt_3649;   // oc8051_tb.v(104)
    output _cvpt_3650;   // oc8051_tb.v(104)
    output _cvpt_3651;   // oc8051_tb.v(104)
    output _cvpt_3652;   // oc8051_tb.v(104)
    output _cvpt_3653;   // oc8051_tb.v(104)
    output _cvpt_3654;   // oc8051_tb.v(104)
    output _cvpt_3655;   // oc8051_tb.v(104)
    output _cvpt_3656;   // oc8051_tb.v(104)
    output _cvpt_3657;   // oc8051_tb.v(104)
    output _cvpt_3658;   // oc8051_tb.v(104)
    output _cvpt_3659;   // oc8051_tb.v(104)
    output _cvpt_3660;   // oc8051_tb.v(104)
    output _cvpt_3661;   // oc8051_tb.v(104)
    output _cvpt_3662;   // oc8051_tb.v(104)
    output _cvpt_3663;   // oc8051_tb.v(104)
    output _cvpt_3664;   // oc8051_tb.v(104)
    output _cvpt_3665;   // oc8051_tb.v(104)
    output _cvpt_3666;   // oc8051_tb.v(104)
    output _cvpt_3667;   // oc8051_tb.v(104)
    output _cvpt_3668;   // oc8051_tb.v(104)
    output _cvpt_3669;   // oc8051_tb.v(104)
    output _cvpt_3670;   // oc8051_tb.v(104)
    output _cvpt_3671;   // oc8051_tb.v(104)
    output _cvpt_3672;   // oc8051_tb.v(104)
    output _cvpt_3673;   // oc8051_tb.v(104)
    output _cvpt_3674;   // oc8051_tb.v(104)
    output _cvpt_3675;   // oc8051_tb.v(104)
    output _cvpt_3676;   // oc8051_tb.v(104)
    output _cvpt_3677;   // oc8051_tb.v(104)
    output _cvpt_3678;   // oc8051_tb.v(104)
    output _cvpt_3679;   // oc8051_tb.v(104)
    output _cvpt_3680;   // oc8051_tb.v(104)
    output _cvpt_3681;   // oc8051_tb.v(104)
    output _cvpt_3682;   // oc8051_tb.v(104)
    output _cvpt_3683;   // oc8051_tb.v(104)
    output _cvpt_3684;   // oc8051_tb.v(104)
    output _cvpt_3685;   // oc8051_tb.v(104)
    output _cvpt_3686;   // oc8051_tb.v(104)
    output _cvpt_3687;   // oc8051_tb.v(104)
    output _cvpt_3688;   // oc8051_tb.v(104)
    output _cvpt_3689;   // oc8051_tb.v(104)
    output _cvpt_3690;   // oc8051_tb.v(104)
    output _cvpt_3691;   // oc8051_tb.v(104)
    output _cvpt_3692;   // oc8051_tb.v(104)
    output _cvpt_3693;   // oc8051_tb.v(104)
    output _cvpt_3694;   // oc8051_tb.v(104)
    output _cvpt_3695;   // oc8051_tb.v(104)
    output _cvpt_3696;   // oc8051_tb.v(104)
    output _cvpt_3697;   // oc8051_tb.v(104)
    output _cvpt_3698;   // oc8051_tb.v(104)
    output _cvpt_3699;   // oc8051_tb.v(104)
    output _cvpt_3700;   // oc8051_tb.v(104)
    output _cvpt_3701;   // oc8051_tb.v(104)
    output _cvpt_3702;   // oc8051_tb.v(104)
    output _cvpt_3703;   // oc8051_tb.v(104)
    output _cvpt_3704;   // oc8051_tb.v(104)
    output _cvpt_3705;   // oc8051_tb.v(104)
    output _cvpt_3706;   // oc8051_tb.v(104)
    output _cvpt_3707;   // oc8051_tb.v(104)
    output _cvpt_3708;   // oc8051_tb.v(104)
    output _cvpt_3709;   // oc8051_tb.v(104)
    output _cvpt_3710;   // oc8051_tb.v(104)
    output _cvpt_3711;   // oc8051_tb.v(104)
    output _cvpt_3712;   // oc8051_tb.v(104)
    output _cvpt_3713;   // oc8051_tb.v(104)
    output _cvpt_3714;   // oc8051_tb.v(104)
    output _cvpt_3715;   // oc8051_tb.v(104)
    output _cvpt_3716;   // oc8051_tb.v(104)
    output _cvpt_3717;   // oc8051_tb.v(104)
    output _cvpt_3718;   // oc8051_tb.v(104)
    output _cvpt_3719;   // oc8051_tb.v(104)
    output _cvpt_3720;   // oc8051_tb.v(104)
    output _cvpt_3721;   // oc8051_tb.v(104)
    output _cvpt_3722;   // oc8051_tb.v(104)
    output _cvpt_3723;   // oc8051_tb.v(104)
    output _cvpt_3724;   // oc8051_tb.v(104)
    output _cvpt_3725;   // oc8051_tb.v(104)
    output _cvpt_3726;   // oc8051_tb.v(104)
    output _cvpt_3727;   // oc8051_tb.v(104)
    output _cvpt_3728;   // oc8051_tb.v(104)
    output _cvpt_3729;   // oc8051_tb.v(104)
    output _cvpt_3730;   // oc8051_tb.v(104)
    output _cvpt_3731;   // oc8051_tb.v(104)
    output _cvpt_3732;   // oc8051_tb.v(104)
    output _cvpt_3733;   // oc8051_tb.v(104)
    output _cvpt_3734;   // oc8051_tb.v(104)
    output _cvpt_3735;   // oc8051_tb.v(104)
    output _cvpt_3736;   // oc8051_tb.v(104)
    output _cvpt_3737;   // oc8051_tb.v(104)
    output _cvpt_3738;   // oc8051_tb.v(104)
    output _cvpt_3739;   // oc8051_tb.v(104)
    output _cvpt_3740;   // oc8051_tb.v(104)
    output _cvpt_3741;   // oc8051_tb.v(104)
    output _cvpt_3742;   // oc8051_tb.v(104)
    output _cvpt_3743;   // oc8051_tb.v(104)
    output _cvpt_3744;   // oc8051_tb.v(104)
    output _cvpt_3745;   // oc8051_tb.v(104)
    output _cvpt_3746;   // oc8051_tb.v(104)
    output _cvpt_3747;   // oc8051_tb.v(104)
    output _cvpt_3748;   // oc8051_tb.v(104)
    output _cvpt_3749;   // oc8051_tb.v(104)
    output _cvpt_3750;   // oc8051_tb.v(104)
    output _cvpt_3751;   // oc8051_tb.v(104)
    output _cvpt_3752;   // oc8051_tb.v(104)
    output _cvpt_3753;   // oc8051_tb.v(104)
    output _cvpt_3754;   // oc8051_tb.v(104)
    output _cvpt_3755;   // oc8051_tb.v(104)
    output _cvpt_3756;   // oc8051_tb.v(104)
    output _cvpt_3757;   // oc8051_tb.v(104)
    output _cvpt_3758;   // oc8051_tb.v(104)
    output _cvpt_3759;   // oc8051_tb.v(104)
    output _cvpt_3760;   // oc8051_tb.v(104)
    output _cvpt_3761;   // oc8051_tb.v(104)
    output _cvpt_3762;   // oc8051_tb.v(104)
    output _cvpt_3763;   // oc8051_tb.v(104)
    output _cvpt_3764;   // oc8051_tb.v(104)
    output _cvpt_3765;   // oc8051_tb.v(104)
    output _cvpt_3766;   // oc8051_tb.v(104)
    output _cvpt_3767;   // oc8051_tb.v(104)
    output _cvpt_3768;   // oc8051_tb.v(104)
    output _cvpt_3769;   // oc8051_tb.v(104)
    output _cvpt_3770;   // oc8051_tb.v(104)
    output _cvpt_3771;   // oc8051_tb.v(104)
    output _cvpt_3772;   // oc8051_tb.v(104)
    output _cvpt_3773;   // oc8051_tb.v(104)
    output _cvpt_3774;   // oc8051_tb.v(104)
    output _cvpt_3775;   // oc8051_tb.v(104)
    output _cvpt_3776;   // oc8051_tb.v(104)
    output _cvpt_3777;   // oc8051_tb.v(104)
    output _cvpt_3778;   // oc8051_tb.v(104)
    output _cvpt_3779;   // oc8051_tb.v(104)
    output _cvpt_3780;   // oc8051_tb.v(104)
    output _cvpt_3781;   // oc8051_tb.v(104)
    output _cvpt_3782;   // oc8051_tb.v(104)
    output _cvpt_3783;   // oc8051_tb.v(104)
    output _cvpt_3784;   // oc8051_tb.v(104)
    output _cvpt_3785;   // oc8051_tb.v(104)
    output _cvpt_3786;   // oc8051_tb.v(104)
    output _cvpt_3787;   // oc8051_tb.v(104)
    output _cvpt_3788;   // oc8051_tb.v(104)
    output _cvpt_3789;   // oc8051_tb.v(104)
    output _cvpt_3790;   // oc8051_tb.v(104)
    output _cvpt_3791;   // oc8051_tb.v(104)
    output _cvpt_3792;   // oc8051_tb.v(104)
    output _cvpt_3793;   // oc8051_tb.v(104)
    output _cvpt_3794;   // oc8051_tb.v(104)
    output _cvpt_3795;   // oc8051_tb.v(104)
    output _cvpt_3796;   // oc8051_tb.v(104)
    output _cvpt_3797;   // oc8051_tb.v(104)
    output _cvpt_3798;   // oc8051_tb.v(104)
    output _cvpt_3799;   // oc8051_tb.v(104)
    output _cvpt_3800;   // oc8051_tb.v(104)
    output _cvpt_3801;   // oc8051_tb.v(104)
    output _cvpt_3802;   // oc8051_tb.v(104)
    output _cvpt_3803;   // oc8051_tb.v(104)
    output _cvpt_3804;   // oc8051_tb.v(104)
    output _cvpt_3805;   // oc8051_tb.v(104)
    output _cvpt_3806;   // oc8051_tb.v(104)
    output _cvpt_3807;   // oc8051_tb.v(104)
    output _cvpt_3808;   // oc8051_tb.v(104)
    output _cvpt_3809;   // oc8051_tb.v(104)
    output _cvpt_3810;   // oc8051_tb.v(104)
    output _cvpt_3811;   // oc8051_tb.v(104)
    output _cvpt_3812;   // oc8051_tb.v(104)
    output _cvpt_3813;   // oc8051_tb.v(104)
    output _cvpt_3814;   // oc8051_tb.v(104)
    output _cvpt_3815;   // oc8051_tb.v(104)
    output _cvpt_3816;   // oc8051_tb.v(104)
    output _cvpt_3817;   // oc8051_tb.v(104)
    output _cvpt_3818;   // oc8051_tb.v(104)
    output _cvpt_3819;   // oc8051_tb.v(104)
    output _cvpt_3820;   // oc8051_tb.v(104)
    output _cvpt_3821;   // oc8051_tb.v(104)
    output _cvpt_3822;   // oc8051_tb.v(104)
    output _cvpt_3823;   // oc8051_tb.v(104)
    output _cvpt_3824;   // oc8051_tb.v(104)
    output _cvpt_3825;   // oc8051_tb.v(104)
    output _cvpt_3826;   // oc8051_tb.v(104)
    output _cvpt_3827;   // oc8051_tb.v(104)
    output _cvpt_3828;   // oc8051_tb.v(104)
    output _cvpt_3829;   // oc8051_tb.v(104)
    output _cvpt_3830;   // oc8051_tb.v(104)
    output _cvpt_3831;   // oc8051_tb.v(104)
    output _cvpt_3832;   // oc8051_tb.v(104)
    output _cvpt_3833;   // oc8051_tb.v(104)
    output _cvpt_3834;   // oc8051_tb.v(104)
    output _cvpt_3835;   // oc8051_tb.v(104)
    output _cvpt_3836;   // oc8051_tb.v(104)
    output _cvpt_3837;   // oc8051_tb.v(104)
    output _cvpt_3838;   // oc8051_tb.v(104)
    output _cvpt_3839;   // oc8051_tb.v(104)
    output _cvpt_3840;   // oc8051_tb.v(104)
    output _cvpt_3841;   // oc8051_tb.v(104)
    output _cvpt_3842;   // oc8051_tb.v(104)
    output _cvpt_3843;   // oc8051_tb.v(104)
    output _cvpt_3844;   // oc8051_tb.v(104)
    output _cvpt_3845;   // oc8051_tb.v(104)
    output _cvpt_3846;   // oc8051_tb.v(104)
    output _cvpt_3847;   // oc8051_tb.v(104)
    output _cvpt_3848;   // oc8051_tb.v(104)
    output _cvpt_3849;   // oc8051_tb.v(104)
    output _cvpt_3850;   // oc8051_tb.v(104)
    output _cvpt_3851;   // oc8051_tb.v(104)
    output _cvpt_3852;   // oc8051_tb.v(104)
    output _cvpt_3853;   // oc8051_tb.v(104)
    output _cvpt_3854;   // oc8051_tb.v(104)
    output _cvpt_3855;   // oc8051_tb.v(104)
    output _cvpt_3856;   // oc8051_tb.v(104)
    output _cvpt_3857;   // oc8051_tb.v(104)
    output _cvpt_3858;   // oc8051_tb.v(104)
    output _cvpt_3859;   // oc8051_tb.v(104)
    output _cvpt_3860;   // oc8051_tb.v(104)
    output _cvpt_3861;   // oc8051_tb.v(104)
    output _cvpt_3862;   // oc8051_tb.v(104)
    output _cvpt_3863;   // oc8051_tb.v(104)
    output _cvpt_3864;   // oc8051_tb.v(104)
    output _cvpt_3865;   // oc8051_tb.v(104)
    output _cvpt_3866;   // oc8051_tb.v(104)
    output _cvpt_3867;   // oc8051_tb.v(104)
    output _cvpt_3868;   // oc8051_tb.v(104)
    output _cvpt_3869;   // oc8051_tb.v(104)
    output _cvpt_3870;   // oc8051_tb.v(104)
    output _cvpt_3871;   // oc8051_tb.v(104)
    output _cvpt_3872;   // oc8051_tb.v(104)
    output _cvpt_3873;   // oc8051_tb.v(104)
    output _cvpt_3874;   // oc8051_tb.v(104)
    output _cvpt_3875;   // oc8051_tb.v(104)
    output _cvpt_3876;   // oc8051_tb.v(104)
    output _cvpt_3877;   // oc8051_tb.v(104)
    output _cvpt_3878;   // oc8051_tb.v(104)
    output _cvpt_3879;   // oc8051_tb.v(104)
    output _cvpt_3880;   // oc8051_tb.v(104)
    output _cvpt_3881;   // oc8051_tb.v(104)
    output _cvpt_3882;   // oc8051_tb.v(104)
    output _cvpt_3883;   // oc8051_tb.v(104)
    output _cvpt_3884;   // oc8051_tb.v(104)
    output _cvpt_3885;   // oc8051_tb.v(104)
    output _cvpt_3886;   // oc8051_tb.v(104)
    output _cvpt_3887;   // oc8051_tb.v(104)
    output _cvpt_3888;   // oc8051_tb.v(104)
    output _cvpt_3889;   // oc8051_tb.v(104)
    output _cvpt_3890;   // oc8051_tb.v(104)
    output _cvpt_3891;   // oc8051_tb.v(104)
    output _cvpt_3892;   // oc8051_tb.v(104)
    output _cvpt_3893;   // oc8051_tb.v(104)
    output _cvpt_3894;   // oc8051_tb.v(104)
    output _cvpt_3895;   // oc8051_tb.v(104)
    output _cvpt_3896;   // oc8051_tb.v(104)
    output _cvpt_3897;   // oc8051_tb.v(104)
    output _cvpt_3898;   // oc8051_tb.v(104)
    output _cvpt_3899;   // oc8051_tb.v(104)
    output _cvpt_3900;   // oc8051_tb.v(104)
    output _cvpt_3901;   // oc8051_tb.v(104)
    output _cvpt_3902;   // oc8051_tb.v(104)
    output _cvpt_3903;   // oc8051_tb.v(104)
    output _cvpt_3904;   // oc8051_tb.v(104)
    output _cvpt_3905;   // oc8051_tb.v(104)
    output _cvpt_3906;   // oc8051_tb.v(104)
    output _cvpt_3907;   // oc8051_tb.v(104)
    output _cvpt_3908;   // oc8051_tb.v(104)
    output _cvpt_3909;   // oc8051_tb.v(104)
    output _cvpt_3910;   // oc8051_tb.v(104)
    output _cvpt_3911;   // oc8051_tb.v(104)
    output _cvpt_3912;   // oc8051_tb.v(104)
    output _cvpt_3913;   // oc8051_tb.v(104)
    output _cvpt_3914;   // oc8051_tb.v(104)
    output _cvpt_3915;   // oc8051_tb.v(104)
    output _cvpt_3916;   // oc8051_tb.v(104)
    output _cvpt_3917;   // oc8051_tb.v(104)
    output _cvpt_3918;   // oc8051_tb.v(104)
    output _cvpt_3919;   // oc8051_tb.v(104)
    output _cvpt_3920;   // oc8051_tb.v(104)
    output _cvpt_3921;   // oc8051_tb.v(104)
    output _cvpt_3922;   // oc8051_tb.v(104)
    output _cvpt_3923;   // oc8051_tb.v(104)
    output _cvpt_3924;   // oc8051_tb.v(104)
    output _cvpt_3925;   // oc8051_tb.v(104)
    output _cvpt_3926;   // oc8051_tb.v(104)
    output _cvpt_3927;   // oc8051_tb.v(104)
    output _cvpt_3928;   // oc8051_tb.v(104)
    output _cvpt_3929;   // oc8051_tb.v(104)
    output _cvpt_3930;   // oc8051_tb.v(104)
    output _cvpt_3931;   // oc8051_tb.v(104)
    output _cvpt_3932;   // oc8051_tb.v(104)
    output _cvpt_3933;   // oc8051_tb.v(104)
    output _cvpt_3934;   // oc8051_tb.v(104)
    output _cvpt_3935;   // oc8051_tb.v(104)
    output _cvpt_3936;   // oc8051_tb.v(104)
    output _cvpt_3937;   // oc8051_tb.v(104)
    output _cvpt_3938;   // oc8051_tb.v(104)
    output _cvpt_3939;   // oc8051_tb.v(104)
    output _cvpt_3940;   // oc8051_tb.v(104)
    output _cvpt_3941;   // oc8051_tb.v(104)
    output _cvpt_3942;   // oc8051_tb.v(104)
    output _cvpt_3943;   // oc8051_tb.v(104)
    output _cvpt_3944;   // oc8051_tb.v(104)
    output _cvpt_3945;   // oc8051_tb.v(104)
    output _cvpt_3946;   // oc8051_tb.v(104)
    output _cvpt_3947;   // oc8051_tb.v(104)
    output _cvpt_3948;   // oc8051_tb.v(104)
    output _cvpt_3949;   // oc8051_tb.v(104)
    output _cvpt_3950;   // oc8051_tb.v(104)
    output _cvpt_3951;   // oc8051_tb.v(104)
    output _cvpt_3952;   // oc8051_tb.v(104)
    output _cvpt_3953;   // oc8051_tb.v(104)
    output _cvpt_3954;   // oc8051_tb.v(104)
    output _cvpt_3955;   // oc8051_tb.v(104)
    output _cvpt_3956;   // oc8051_tb.v(104)
    output _cvpt_3957;   // oc8051_tb.v(104)
    output _cvpt_3958;   // oc8051_tb.v(104)
    output _cvpt_3959;   // oc8051_tb.v(104)
    output _cvpt_3960;   // oc8051_tb.v(104)
    output _cvpt_3961;   // oc8051_tb.v(104)
    output _cvpt_3962;   // oc8051_tb.v(104)
    output _cvpt_3963;   // oc8051_tb.v(104)
    output _cvpt_3964;   // oc8051_tb.v(104)
    output _cvpt_3965;   // oc8051_tb.v(104)
    output _cvpt_3966;   // oc8051_tb.v(104)
    output _cvpt_3967;   // oc8051_tb.v(104)
    output _cvpt_3968;   // oc8051_tb.v(104)
    output _cvpt_3969;   // oc8051_tb.v(104)
    output _cvpt_3970;   // oc8051_tb.v(104)
    output _cvpt_3971;   // oc8051_tb.v(104)
    output _cvpt_3972;   // oc8051_tb.v(104)
    output _cvpt_3973;   // oc8051_tb.v(104)
    output _cvpt_3974;   // oc8051_tb.v(104)
    output _cvpt_3975;   // oc8051_tb.v(104)
    output _cvpt_3976;   // oc8051_tb.v(104)
    output _cvpt_3977;   // oc8051_tb.v(104)
    output _cvpt_3978;   // oc8051_tb.v(104)
    output _cvpt_3979;   // oc8051_tb.v(104)
    output _cvpt_3980;   // oc8051_tb.v(104)
    output _cvpt_3981;   // oc8051_tb.v(104)
    output _cvpt_3982;   // oc8051_tb.v(104)
    output _cvpt_3983;   // oc8051_tb.v(104)
    output _cvpt_3984;   // oc8051_tb.v(104)
    output _cvpt_3985;   // oc8051_tb.v(104)
    output _cvpt_3986;   // oc8051_tb.v(104)
    output _cvpt_3987;   // oc8051_tb.v(104)
    output _cvpt_3988;   // oc8051_tb.v(104)
    output _cvpt_3989;   // oc8051_tb.v(104)
    output _cvpt_3990;   // oc8051_tb.v(104)
    output _cvpt_3991;   // oc8051_tb.v(104)
    output _cvpt_3992;   // oc8051_tb.v(104)
    output _cvpt_3993;   // oc8051_tb.v(104)
    output _cvpt_3994;   // oc8051_tb.v(104)
    output _cvpt_3995;   // oc8051_tb.v(104)
    output _cvpt_3996;   // oc8051_tb.v(104)
    output _cvpt_3997;   // oc8051_tb.v(104)
    output _cvpt_3998;   // oc8051_tb.v(104)
    output _cvpt_3999;   // oc8051_tb.v(104)
    output _cvpt_4000;   // oc8051_tb.v(104)
    output _cvpt_4001;   // oc8051_tb.v(104)
    output _cvpt_4002;   // oc8051_tb.v(104)
    output _cvpt_4003;   // oc8051_tb.v(104)
    output _cvpt_4004;   // oc8051_tb.v(104)
    output _cvpt_4005;   // oc8051_tb.v(104)
    output _cvpt_4006;   // oc8051_tb.v(104)
    output _cvpt_4007;   // oc8051_tb.v(104)
    output _cvpt_4008;   // oc8051_tb.v(104)
    output _cvpt_4009;   // oc8051_tb.v(104)
    output _cvpt_4010;   // oc8051_tb.v(104)
    output _cvpt_4011;   // oc8051_tb.v(104)
    output _cvpt_4012;   // oc8051_tb.v(104)
    output _cvpt_4013;   // oc8051_tb.v(104)
    output _cvpt_4014;   // oc8051_tb.v(104)
    output _cvpt_4015;   // oc8051_tb.v(104)
    output _cvpt_4016;   // oc8051_tb.v(104)
    output _cvpt_4017;   // oc8051_tb.v(104)
    output _cvpt_4018;   // oc8051_tb.v(104)
    output _cvpt_4019;   // oc8051_tb.v(104)
    output _cvpt_4020;   // oc8051_tb.v(104)
    output _cvpt_4021;   // oc8051_tb.v(104)
    output _cvpt_4022;   // oc8051_tb.v(104)
    output _cvpt_4023;   // oc8051_tb.v(104)
    output _cvpt_4024;   // oc8051_tb.v(104)
    output _cvpt_4025;   // oc8051_tb.v(104)
    output _cvpt_4026;   // oc8051_tb.v(104)
    output _cvpt_4027;   // oc8051_tb.v(104)
    output _cvpt_4028;   // oc8051_tb.v(104)
    output _cvpt_4029;   // oc8051_tb.v(104)
    output _cvpt_4030;   // oc8051_tb.v(104)
    output _cvpt_4031;   // oc8051_tb.v(104)
    output _cvpt_4032;   // oc8051_tb.v(104)
    output _cvpt_4033;   // oc8051_tb.v(104)
    output _cvpt_4034;   // oc8051_tb.v(104)
    output _cvpt_4035;   // oc8051_tb.v(104)
    output _cvpt_4036;   // oc8051_tb.v(104)
    output _cvpt_4037;   // oc8051_tb.v(104)
    output _cvpt_4038;   // oc8051_tb.v(104)
    output _cvpt_4039;   // oc8051_tb.v(104)
    output _cvpt_4040;   // oc8051_tb.v(104)
    output _cvpt_4041;   // oc8051_tb.v(104)
    output _cvpt_4042;   // oc8051_tb.v(104)
    output _cvpt_4043;   // oc8051_tb.v(104)
    output _cvpt_4044;   // oc8051_tb.v(104)
    output _cvpt_4045;   // oc8051_tb.v(104)
    output _cvpt_4046;   // oc8051_tb.v(104)
    output _cvpt_4047;   // oc8051_tb.v(104)
    output _cvpt_4048;   // oc8051_tb.v(104)
    output _cvpt_4049;   // oc8051_tb.v(104)
    output _cvpt_4050;   // oc8051_tb.v(104)
    output _cvpt_4051;   // oc8051_tb.v(104)
    output _cvpt_4052;   // oc8051_tb.v(104)
    output _cvpt_4053;   // oc8051_tb.v(104)
    output _cvpt_4054;   // oc8051_tb.v(104)
    output _cvpt_4055;   // oc8051_tb.v(104)
    output _cvpt_4056;   // oc8051_tb.v(104)
    output _cvpt_4057;   // oc8051_tb.v(104)
    output _cvpt_4058;   // oc8051_tb.v(104)
    output _cvpt_4059;   // oc8051_tb.v(104)
    output _cvpt_4060;   // oc8051_tb.v(104)
    output _cvpt_4061;   // oc8051_tb.v(104)
    output _cvpt_4062;   // oc8051_tb.v(104)
    output _cvpt_4063;   // oc8051_tb.v(104)
    output _cvpt_4064;   // oc8051_tb.v(104)
    output _cvpt_4065;   // oc8051_tb.v(104)
    output _cvpt_4066;   // oc8051_tb.v(104)
    output _cvpt_4067;   // oc8051_tb.v(104)
    output _cvpt_4068;   // oc8051_tb.v(104)
    output _cvpt_4069;   // oc8051_tb.v(104)
    output _cvpt_4070;   // oc8051_tb.v(104)
    output _cvpt_4071;   // oc8051_tb.v(104)
    output _cvpt_4072;   // oc8051_tb.v(104)
    output _cvpt_4073;   // oc8051_tb.v(104)
    output _cvpt_4074;   // oc8051_tb.v(104)
    output _cvpt_4075;   // oc8051_tb.v(104)
    output _cvpt_4076;   // oc8051_tb.v(104)
    output _cvpt_4077;   // oc8051_tb.v(104)
    output _cvpt_4078;   // oc8051_tb.v(104)
    output _cvpt_4079;   // oc8051_tb.v(104)
    output _cvpt_4080;   // oc8051_tb.v(104)
    output _cvpt_4081;   // oc8051_tb.v(104)
    output _cvpt_4082;   // oc8051_tb.v(104)
    output _cvpt_4083;   // oc8051_tb.v(104)
    output _cvpt_4084;   // oc8051_tb.v(104)
    output _cvpt_4085;   // oc8051_tb.v(104)
    output _cvpt_4086;   // oc8051_tb.v(104)
    output _cvpt_4087;   // oc8051_tb.v(104)
    output _cvpt_4088;   // oc8051_tb.v(104)
    output _cvpt_4089;   // oc8051_tb.v(104)
    output _cvpt_4090;   // oc8051_tb.v(104)
    output _cvpt_4091;   // oc8051_tb.v(104)
    output _cvpt_4092;   // oc8051_tb.v(104)
    output _cvpt_4093;   // oc8051_tb.v(104)
    output _cvpt_4094;   // oc8051_tb.v(104)
    output _cvpt_4095;   // oc8051_tb.v(104)
    output _cvpt_4096;   // oc8051_tb.v(104)
    output _cvpt_4097;   // oc8051_tb.v(104)
    output _cvpt_4098;   // oc8051_tb.v(104)
    output _cvpt_4099;   // oc8051_tb.v(104)
    output _cvpt_4100;   // oc8051_tb.v(104)
    output _cvpt_4101;   // oc8051_tb.v(104)
    output _cvpt_4102;   // oc8051_tb.v(104)
    output _cvpt_4103;   // oc8051_tb.v(104)
    output _cvpt_4104;   // oc8051_tb.v(104)
    output _cvpt_4105;   // oc8051_tb.v(104)
    output _cvpt_4106;   // oc8051_tb.v(104)
    output _cvpt_4107;   // oc8051_tb.v(104)
    output _cvpt_4108;   // oc8051_tb.v(104)
    output _cvpt_4109;   // oc8051_tb.v(104)
    output _cvpt_4110;   // oc8051_tb.v(104)
    output _cvpt_4111;   // oc8051_tb.v(104)
    output _cvpt_4112;   // oc8051_tb.v(104)
    output _cvpt_4113;   // oc8051_tb.v(104)
    output _cvpt_4114;   // oc8051_tb.v(104)
    output _cvpt_4115;   // oc8051_tb.v(104)
    output _cvpt_4116;   // oc8051_tb.v(104)
    output _cvpt_4117;   // oc8051_tb.v(104)
    output _cvpt_4118;   // oc8051_tb.v(104)
    output _cvpt_4119;   // oc8051_tb.v(104)
    output _cvpt_4120;   // oc8051_tb.v(104)
    output _cvpt_4121;   // oc8051_tb.v(104)
    output _cvpt_4122;   // oc8051_tb.v(104)
    output _cvpt_4123;   // oc8051_tb.v(104)
    output _cvpt_4124;   // oc8051_tb.v(104)
    output _cvpt_4125;   // oc8051_tb.v(104)
    output _cvpt_4126;   // oc8051_tb.v(104)
    output _cvpt_4127;   // oc8051_tb.v(104)
    output _cvpt_4128;   // oc8051_tb.v(104)
    output _cvpt_4129;   // oc8051_tb.v(104)
    output _cvpt_4130;   // oc8051_tb.v(104)
    output _cvpt_4131;   // oc8051_tb.v(104)
    output _cvpt_4132;   // oc8051_tb.v(104)
    output _cvpt_4133;   // oc8051_tb.v(104)
    output _cvpt_4134;   // oc8051_tb.v(104)
    output _cvpt_4135;   // oc8051_tb.v(104)
    output _cvpt_4136;   // oc8051_tb.v(104)
    output _cvpt_4137;   // oc8051_tb.v(104)
    output _cvpt_4138;   // oc8051_tb.v(104)
    output _cvpt_4139;   // oc8051_tb.v(104)
    output _cvpt_4140;   // oc8051_tb.v(104)
    output _cvpt_4141;   // oc8051_tb.v(104)
    output _cvpt_4142;   // oc8051_tb.v(104)
    output _cvpt_4143;   // oc8051_tb.v(104)
    output _cvpt_4144;   // oc8051_tb.v(104)
    output _cvpt_4145;   // oc8051_tb.v(104)
    output _cvpt_4146;   // oc8051_tb.v(104)
    output _cvpt_4147;   // oc8051_tb.v(104)
    output _cvpt_4148;   // oc8051_tb.v(104)
    output _cvpt_4149;   // oc8051_tb.v(104)
    output _cvpt_4150;   // oc8051_tb.v(104)
    output _cvpt_4151;   // oc8051_tb.v(104)
    output _cvpt_4152;   // oc8051_tb.v(104)
    output _cvpt_4153;   // oc8051_tb.v(104)
    output _cvpt_4154;   // oc8051_tb.v(104)
    output _cvpt_4155;   // oc8051_tb.v(104)
    output _cvpt_4156;   // oc8051_tb.v(104)
    output _cvpt_4157;   // oc8051_tb.v(104)
    output _cvpt_4158;   // oc8051_tb.v(104)
    output _cvpt_4159;   // oc8051_tb.v(104)
    output _cvpt_4160;   // oc8051_tb.v(104)
    output _cvpt_4161;   // oc8051_tb.v(104)
    output _cvpt_4162;   // oc8051_tb.v(104)
    output _cvpt_4163;   // oc8051_tb.v(104)
    output _cvpt_4164;   // oc8051_tb.v(104)
    output _cvpt_4165;   // oc8051_tb.v(104)
    output _cvpt_4166;   // oc8051_tb.v(104)
    output _cvpt_4167;   // oc8051_tb.v(104)
    output _cvpt_4168;   // oc8051_tb.v(104)
    output _cvpt_4169;   // oc8051_tb.v(104)
    output _cvpt_4170;   // oc8051_tb.v(104)
    output _cvpt_4171;   // oc8051_tb.v(104)
    output _cvpt_4172;   // oc8051_tb.v(104)
    output _cvpt_4173;   // oc8051_tb.v(104)
    output _cvpt_4174;   // oc8051_tb.v(104)
    output _cvpt_4175;   // oc8051_tb.v(104)
    output _cvpt_4176;   // oc8051_tb.v(104)
    output _cvpt_4177;   // oc8051_tb.v(104)
    output _cvpt_4178;   // oc8051_tb.v(104)
    output _cvpt_4179;   // oc8051_tb.v(104)
    output _cvpt_4180;   // oc8051_tb.v(104)
    output _cvpt_4181;   // oc8051_tb.v(104)
    output _cvpt_4182;   // oc8051_tb.v(104)
    output _cvpt_4183;   // oc8051_tb.v(104)
    output _cvpt_4184;   // oc8051_tb.v(104)
    output _cvpt_4185;   // oc8051_tb.v(104)
    output _cvpt_4186;   // oc8051_tb.v(104)
    output _cvpt_4187;   // oc8051_tb.v(104)
    output _cvpt_4188;   // oc8051_tb.v(104)
    output _cvpt_4189;   // oc8051_tb.v(104)
    output _cvpt_4190;   // oc8051_tb.v(104)
    output _cvpt_4191;   // oc8051_tb.v(104)
    output _cvpt_4192;   // oc8051_tb.v(104)
    output _cvpt_4193;   // oc8051_tb.v(104)
    output _cvpt_4194;   // oc8051_tb.v(104)
    output _cvpt_4195;   // oc8051_tb.v(104)
    output _cvpt_4196;   // oc8051_tb.v(104)
    output _cvpt_4197;   // oc8051_tb.v(104)
    output _cvpt_4198;   // oc8051_tb.v(104)
    output _cvpt_4199;   // oc8051_tb.v(104)
    output _cvpt_4200;   // oc8051_tb.v(104)
    output _cvpt_4201;   // oc8051_tb.v(104)
    output _cvpt_4202;   // oc8051_tb.v(104)
    output _cvpt_4203;   // oc8051_tb.v(104)
    output _cvpt_4204;   // oc8051_tb.v(104)
    output _cvpt_4205;   // oc8051_tb.v(104)
    output _cvpt_4206;   // oc8051_tb.v(104)
    output _cvpt_4207;   // oc8051_tb.v(104)
    output _cvpt_4208;   // oc8051_tb.v(104)
    output _cvpt_4209;   // oc8051_tb.v(104)
    output _cvpt_4210;   // oc8051_tb.v(104)
    output _cvpt_4211;   // oc8051_tb.v(104)
    output _cvpt_4212;   // oc8051_tb.v(104)
    output _cvpt_4213;   // oc8051_tb.v(104)
    output _cvpt_4214;   // oc8051_tb.v(104)
    output _cvpt_4215;   // oc8051_tb.v(104)
    output _cvpt_4216;   // oc8051_tb.v(104)
    output _cvpt_4217;   // oc8051_tb.v(104)
    output _cvpt_4218;   // oc8051_tb.v(104)
    output _cvpt_4219;   // oc8051_tb.v(104)
    output _cvpt_4220;   // oc8051_tb.v(104)
    output _cvpt_4221;   // oc8051_tb.v(104)
    output _cvpt_4222;   // oc8051_tb.v(104)
    output _cvpt_4223;   // oc8051_tb.v(104)
    output _cvpt_4224;   // oc8051_tb.v(104)
    output _cvpt_4225;   // oc8051_tb.v(104)
    output _cvpt_4226;   // oc8051_tb.v(104)
    output _cvpt_4227;   // oc8051_tb.v(104)
    output _cvpt_4228;   // oc8051_tb.v(104)
    output _cvpt_4229;   // oc8051_tb.v(104)
    output _cvpt_4230;   // oc8051_tb.v(104)
    output _cvpt_4231;   // oc8051_tb.v(104)
    output _cvpt_4232;   // oc8051_tb.v(104)
    output _cvpt_4233;   // oc8051_tb.v(104)
    output _cvpt_4234;   // oc8051_tb.v(104)
    output _cvpt_4235;   // oc8051_tb.v(104)
    output _cvpt_4236;   // oc8051_tb.v(104)
    output _cvpt_4237;   // oc8051_tb.v(104)
    output _cvpt_4238;   // oc8051_tb.v(104)
    output _cvpt_4239;   // oc8051_tb.v(104)
    output _cvpt_4240;   // oc8051_tb.v(104)
    output _cvpt_4241;   // oc8051_tb.v(104)
    output _cvpt_4242;   // oc8051_tb.v(104)
    output _cvpt_4243;   // oc8051_tb.v(104)
    output _cvpt_4244;   // oc8051_tb.v(104)
    output _cvpt_4245;   // oc8051_tb.v(104)
    output _cvpt_4246;   // oc8051_tb.v(104)
    output _cvpt_4247;   // oc8051_tb.v(104)
    output _cvpt_4248;   // oc8051_tb.v(104)
    output _cvpt_4249;   // oc8051_tb.v(104)
    output _cvpt_4250;   // oc8051_tb.v(104)
    output _cvpt_4251;   // oc8051_tb.v(104)
    output _cvpt_4252;   // oc8051_tb.v(104)
    output _cvpt_4253;   // oc8051_tb.v(104)
    output _cvpt_4254;   // oc8051_tb.v(104)
    output _cvpt_4255;   // oc8051_tb.v(104)
    output _cvpt_4256;   // oc8051_tb.v(104)
    output _cvpt_4257;   // oc8051_tb.v(104)
    output _cvpt_4258;   // oc8051_tb.v(104)
    output _cvpt_4259;   // oc8051_tb.v(104)
    output _cvpt_4260;   // oc8051_tb.v(104)
    output _cvpt_4261;   // oc8051_tb.v(104)
    output _cvpt_4262;   // oc8051_tb.v(104)
    output _cvpt_4263;   // oc8051_tb.v(104)
    output _cvpt_4264;   // oc8051_tb.v(104)
    output _cvpt_4265;   // oc8051_tb.v(104)
    output _cvpt_4266;   // oc8051_tb.v(104)
    output _cvpt_4267;   // oc8051_tb.v(104)
    output _cvpt_4268;   // oc8051_tb.v(104)
    output _cvpt_4269;   // oc8051_tb.v(104)
    output _cvpt_4270;   // oc8051_tb.v(104)
    output _cvpt_4271;   // oc8051_tb.v(104)
    output _cvpt_4272;   // oc8051_tb.v(104)
    output _cvpt_4273;   // oc8051_tb.v(104)
    output _cvpt_4274;   // oc8051_tb.v(104)
    output _cvpt_4275;   // oc8051_tb.v(104)
    output _cvpt_4276;   // oc8051_tb.v(104)
    output _cvpt_4277;   // oc8051_tb.v(104)
    output _cvpt_4278;   // oc8051_tb.v(104)
    output _cvpt_4279;   // oc8051_tb.v(104)
    output _cvpt_4280;   // oc8051_tb.v(104)
    output _cvpt_4281;   // oc8051_tb.v(104)
    output _cvpt_4282;   // oc8051_tb.v(104)
    output _cvpt_4283;   // oc8051_tb.v(104)
    output _cvpt_4284;   // oc8051_tb.v(104)
    output _cvpt_4285;   // oc8051_tb.v(104)
    output _cvpt_4286;   // oc8051_tb.v(104)
    output _cvpt_4287;   // oc8051_tb.v(104)
    output _cvpt_4288;   // oc8051_tb.v(104)
    output _cvpt_4289;   // oc8051_tb.v(104)
    output _cvpt_4290;   // oc8051_tb.v(104)
    output _cvpt_4291;   // oc8051_tb.v(104)
    output _cvpt_4292;   // oc8051_tb.v(104)
    output _cvpt_4293;   // oc8051_tb.v(104)
    output _cvpt_4294;   // oc8051_tb.v(104)
    output _cvpt_4295;   // oc8051_tb.v(104)
    output _cvpt_4296;   // oc8051_tb.v(104)
    output _cvpt_4297;   // oc8051_tb.v(104)
    output _cvpt_4298;   // oc8051_tb.v(104)
    output _cvpt_4299;   // oc8051_tb.v(104)
    output _cvpt_4300;   // oc8051_tb.v(104)
    output _cvpt_4301;   // oc8051_tb.v(104)
    output _cvpt_4302;   // oc8051_tb.v(104)
    output _cvpt_4303;   // oc8051_tb.v(104)
    output _cvpt_4304;   // oc8051_tb.v(104)
    output _cvpt_4305;   // oc8051_tb.v(104)
    output _cvpt_4306;   // oc8051_tb.v(104)
    output _cvpt_4307;   // oc8051_tb.v(104)
    output _cvpt_4308;   // oc8051_tb.v(104)
    output _cvpt_4309;   // oc8051_tb.v(104)
    output _cvpt_4310;   // oc8051_tb.v(104)
    output _cvpt_4311;   // oc8051_tb.v(104)
    output _cvpt_4312;   // oc8051_tb.v(104)
    output _cvpt_4313;   // oc8051_tb.v(104)
    output _cvpt_4314;   // oc8051_tb.v(104)
    output _cvpt_4315;   // oc8051_tb.v(104)
    output _cvpt_4316;   // oc8051_tb.v(104)
    output _cvpt_4317;   // oc8051_tb.v(104)
    output _cvpt_4318;   // oc8051_tb.v(104)
    output _cvpt_4319;   // oc8051_tb.v(104)
    output _cvpt_4320;   // oc8051_tb.v(104)
    output _cvpt_4321;   // oc8051_tb.v(104)
    output _cvpt_4322;   // oc8051_tb.v(104)
    output _cvpt_4323;   // oc8051_tb.v(104)
    output _cvpt_4324;   // oc8051_tb.v(104)
    output _cvpt_4325;   // oc8051_tb.v(104)
    output _cvpt_4326;   // oc8051_tb.v(104)
    output _cvpt_4327;   // oc8051_tb.v(104)
    output _cvpt_4328;   // oc8051_tb.v(104)
    output _cvpt_4329;   // oc8051_tb.v(104)
    output _cvpt_4330;   // oc8051_tb.v(104)
    output _cvpt_4331;   // oc8051_tb.v(104)
    output _cvpt_4332;   // oc8051_tb.v(104)
    output _cvpt_4333;   // oc8051_tb.v(104)
    output _cvpt_4334;   // oc8051_tb.v(104)
    output _cvpt_4335;   // oc8051_tb.v(104)
    output _cvpt_4336;   // oc8051_tb.v(104)
    output _cvpt_4337;   // oc8051_tb.v(104)
    output _cvpt_4338;   // oc8051_tb.v(104)
    output _cvpt_4339;   // oc8051_tb.v(104)
    output _cvpt_4340;   // oc8051_tb.v(104)
    output _cvpt_4341;   // oc8051_tb.v(104)
    output _cvpt_4342;   // oc8051_tb.v(104)
    output _cvpt_4343;   // oc8051_tb.v(104)
    output _cvpt_4344;   // oc8051_tb.v(104)
    output _cvpt_4345;   // oc8051_tb.v(104)
    output _cvpt_4346;   // oc8051_tb.v(104)
    output _cvpt_4347;   // oc8051_tb.v(104)
    output _cvpt_4348;   // oc8051_tb.v(104)
    output _cvpt_4349;   // oc8051_tb.v(104)
    output _cvpt_4350;   // oc8051_tb.v(104)
    output _cvpt_4351;   // oc8051_tb.v(104)
    output _cvpt_4352;   // oc8051_tb.v(104)
    output _cvpt_4353;   // oc8051_tb.v(104)
    output _cvpt_4354;   // oc8051_tb.v(104)
    output _cvpt_4355;   // oc8051_tb.v(104)
    output _cvpt_4356;   // oc8051_tb.v(104)
    output _cvpt_4357;   // oc8051_tb.v(104)
    output _cvpt_4358;   // oc8051_tb.v(104)
    output _cvpt_4359;   // oc8051_tb.v(104)
    output _cvpt_4360;   // oc8051_tb.v(104)
    output _cvpt_4361;   // oc8051_tb.v(104)
    output _cvpt_4362;   // oc8051_tb.v(104)
    output _cvpt_4363;   // oc8051_tb.v(104)
    output _cvpt_4364;   // oc8051_tb.v(104)
    output _cvpt_4365;   // oc8051_tb.v(104)
    output _cvpt_4366;   // oc8051_tb.v(104)
    output _cvpt_4367;   // oc8051_tb.v(104)
    output _cvpt_4368;   // oc8051_tb.v(104)
    output _cvpt_4369;   // oc8051_tb.v(104)
    output _cvpt_4370;   // oc8051_tb.v(104)
    output _cvpt_4371;   // oc8051_tb.v(104)
    output _cvpt_4372;   // oc8051_tb.v(104)
    output _cvpt_4373;   // oc8051_tb.v(104)
    output _cvpt_4374;   // oc8051_tb.v(104)
    output _cvpt_4375;   // oc8051_tb.v(104)
    output _cvpt_4376;   // oc8051_tb.v(104)
    output _cvpt_4377;   // oc8051_tb.v(104)
    output _cvpt_4378;   // oc8051_tb.v(104)
    output _cvpt_4379;   // oc8051_tb.v(104)
    output _cvpt_4380;   // oc8051_tb.v(104)
    output _cvpt_4381;   // oc8051_tb.v(104)
    output _cvpt_4382;   // oc8051_tb.v(104)
    output _cvpt_4383;   // oc8051_tb.v(104)
    output _cvpt_4384;   // oc8051_tb.v(104)
    output _cvpt_4385;   // oc8051_tb.v(104)
    output _cvpt_4386;   // oc8051_tb.v(104)
    output _cvpt_4387;   // oc8051_tb.v(104)
    output _cvpt_4388;   // oc8051_tb.v(104)
    output _cvpt_4389;   // oc8051_tb.v(104)
    output _cvpt_4390;   // oc8051_tb.v(104)
    output _cvpt_4391;   // oc8051_tb.v(104)
    output _cvpt_4392;   // oc8051_tb.v(104)
    output _cvpt_4393;   // oc8051_tb.v(104)
    output _cvpt_4394;   // oc8051_tb.v(104)
    output _cvpt_4395;   // oc8051_tb.v(104)
    output _cvpt_4396;   // oc8051_tb.v(104)
    output _cvpt_4397;   // oc8051_tb.v(104)
    output _cvpt_4398;   // oc8051_tb.v(104)
    output _cvpt_4399;   // oc8051_tb.v(104)
    output _cvpt_4400;   // oc8051_tb.v(104)
    output _cvpt_4401;   // oc8051_tb.v(104)
    output _cvpt_4402;   // oc8051_tb.v(104)
    output _cvpt_4403;   // oc8051_tb.v(104)
    output _cvpt_4404;   // oc8051_tb.v(104)
    output _cvpt_4405;   // oc8051_tb.v(104)
    output _cvpt_4406;   // oc8051_tb.v(104)
    output _cvpt_4407;   // oc8051_tb.v(104)
    output _cvpt_4408;   // oc8051_tb.v(104)
    output _cvpt_4409;   // oc8051_tb.v(104)
    output _cvpt_4410;   // oc8051_tb.v(104)
    output _cvpt_4411;   // oc8051_tb.v(104)
    output _cvpt_4412;   // oc8051_tb.v(104)
    output _cvpt_4413;   // oc8051_tb.v(104)
    output _cvpt_4414;   // oc8051_tb.v(104)
    output _cvpt_4415;   // oc8051_tb.v(104)
    output _cvpt_4416;   // oc8051_tb.v(104)
    output _cvpt_4417;   // oc8051_tb.v(104)
    output _cvpt_4418;   // oc8051_tb.v(104)
    output _cvpt_4419;   // oc8051_tb.v(104)
    output _cvpt_4420;   // oc8051_tb.v(104)
    output _cvpt_4421;   // oc8051_tb.v(104)
    output _cvpt_4422;   // oc8051_tb.v(104)
    output _cvpt_4423;   // oc8051_tb.v(104)
    output _cvpt_4424;   // oc8051_tb.v(104)
    output _cvpt_4425;   // oc8051_tb.v(104)
    output _cvpt_4426;   // oc8051_tb.v(104)
    output _cvpt_4427;   // oc8051_tb.v(104)
    output _cvpt_4428;   // oc8051_tb.v(104)
    output _cvpt_4429;   // oc8051_tb.v(104)
    output _cvpt_4430;   // oc8051_tb.v(104)
    output _cvpt_4431;   // oc8051_tb.v(104)
    output _cvpt_4432;   // oc8051_tb.v(104)
    output _cvpt_4433;   // oc8051_tb.v(104)
    output _cvpt_4434;   // oc8051_tb.v(104)
    output _cvpt_4435;   // oc8051_tb.v(104)
    output _cvpt_4436;   // oc8051_tb.v(104)
    
    wire [2047:0]\oc8051_xiommu1/exp_exp ;   // oc8051_xiommu.v(67)
    wire [7:0]p0_in;   // oc8051_tb.v(113)
    wire [7:0]p1_in;   // oc8051_tb.v(113)
    wire [7:0]p2_in;   // oc8051_tb.v(113)
    wire [15:0]ext_addr;   // oc8051_tb.v(114)
    wire write;   // oc8051_tb.v(115)
    wire write_xram;   // oc8051_tb.v(115)
    wire write_uart;   // oc8051_tb.v(115)
    wire txd;   // oc8051_tb.v(115)
    wire int0;   // oc8051_tb.v(115)
    wire int1;   // oc8051_tb.v(115)
    wire stb_o;   // oc8051_tb.v(115)
    wire ack_i;   // oc8051_tb.v(115)
    wire ack_xram;   // oc8051_tb.v(116)
    wire ack_uart;   // oc8051_tb.v(116)
    wire iack_i;   // oc8051_tb.v(116)
    wire [7:0]data_in;   // oc8051_tb.v(117)
    wire [7:0]data_out;   // oc8051_tb.v(117)
    wire [7:0]p0_out;   // oc8051_tb.v(117)
    wire [7:0]p1_out;   // oc8051_tb.v(117)
    wire [7:0]p2_out;   // oc8051_tb.v(117)
    wire [7:0]p3_out;   // oc8051_tb.v(117)
    wire [7:0]data_out_uart;   // oc8051_tb.v(117)
    wire [7:0]data_out_xram;   // oc8051_tb.v(117)
    wire [7:0]p3_in;   // oc8051_tb.v(117)
    wire priv_lvl;   // oc8051_tb.v(119)
    wire [15:0]dpc_ot;   // oc8051_tb.v(120)
    wire [31:0]idat_i;   // oc8051_tb.v(125)
    wire [2047:0]\oc8051_xiommu1/exp_m ;   // oc8051_xiommu.v(67)
    wire [127:0]\oc8051_xiommu1/aes_key1 ;   // oc8051_xiommu.v(66)
    wire [127:0]\oc8051_xiommu1/aes_key0 ;   // oc8051_xiommu.v(66)
    wire [127:0]\oc8051_xiommu1/aes_ctr ;   // oc8051_xiommu.v(66)
    wire [15:0]\oc8051_xiommu1/memwr_len ;   // oc8051_xiommu.v(80)
    wire [15:0]\oc8051_xiommu1/memwr_wraddr ;   // oc8051_xiommu.v(80)
    wire [15:0]\oc8051_xiommu1/memwr_rdaddr ;   // oc8051_xiommu.v(80)
    wire [15:0]\oc8051_xiommu1/exp_addr ;   // oc8051_xiommu.v(65)
    wire [15:0]\oc8051_xiommu1/sha_len ;   // oc8051_xiommu.v(65)
    wire [15:0]\oc8051_xiommu1/sha_wraddr ;   // oc8051_xiommu.v(65)
    wire [15:0]\oc8051_xiommu1/sha_rdaddr ;   // oc8051_xiommu.v(65)
    wire [15:0]\oc8051_xiommu1/aes_len ;   // oc8051_xiommu.v(65)
    wire [15:0]\oc8051_xiommu1/aes_addr ;   // oc8051_xiommu.v(65)
    wire \oc8051_xiommu1/memwr_step ;   // oc8051_xiommu.v(79)
    wire \oc8051_xiommu1/exp_step ;   // oc8051_xiommu.v(64)
    wire \oc8051_xiommu1/sha_step ;   // oc8051_xiommu.v(64)
    wire \oc8051_xiommu1/aes_step ;   // oc8051_xiommu.v(64)
    wire [1:0]\oc8051_xiommu1/memwr_state ;   // oc8051_xiommu.v(78)
    wire [1:0]\oc8051_xiommu1/exp_state ;   // oc8051_xiommu.v(63)
    wire [2:0]\oc8051_xiommu1/sha_state ;   // oc8051_xiommu.v(62)
    wire [1:0]\oc8051_xiommu1/aes_state ;   // oc8051_xiommu.v(61)
    wire \oc8051_xiommu1/ack_ia ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/ack_pt ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/ia_addr_range ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/pt_addr_range ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/priv_lvl ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/rd_en ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/wr_en ;   // oc8051_xiommu.v(73)
    wire \oc8051_xiommu1/memwr_addr_range ;   // oc8051_xiommu.v(72)
    wire \oc8051_xiommu1/exp_addr_range ;   // oc8051_xiommu.v(72)
    wire \oc8051_xiommu1/sha_addr_range ;   // oc8051_xiommu.v(72)
    wire \oc8051_xiommu1/aes_addr_range ;   // oc8051_xiommu.v(72)
    wire \oc8051_xiommu1/proc0_stb_xram ;   // oc8051_xiommu.v(71)
    wire \oc8051_xiommu1/proc1_stb_xram ;   // oc8051_xiommu.v(71)
    wire \oc8051_xiommu1/ack_memwr ;   // oc8051_xiommu.v(70)
    wire \oc8051_xiommu1/ack_exp ;   // oc8051_xiommu.v(70)
    wire \oc8051_xiommu1/ack_sha ;   // oc8051_xiommu.v(70)
    wire \oc8051_xiommu1/ack_aes ;   // oc8051_xiommu.v(70)
    wire \oc8051_xiommu1/write_pt ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write_memwr ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write_exp ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write_sha ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write_aes ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write0_xram ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/write1_xram ;   // oc8051_xiommu.v(69)
    wire \oc8051_xiommu1/exp_valid ;   // oc8051_xiommu.v(64)
    wire \oc8051_xiommu1/sha_core_assumps_valid ;   // oc8051_xiommu.v(64)
    wire \oc8051_top_1/oc8051_decoder1/stb_i ;   // oc8051_decoder.v(166)
    wire [2:0]\oc8051_top_1/oc8051_decoder1/ram_rd_sel_r ;   // oc8051_decoder.v(164)
    wire [7:0]\oc8051_top_1/oc8051_decoder1/op ;   // oc8051_decoder.v(162)
    wire [2:0]\oc8051_top_1/oc8051_decoder1/ram_rd_sel ;   // oc8051_decoder.v(154)
    wire [2:0]\oc8051_top_1/oc8051_decoder1/ram_wr_sel ;   // oc8051_decoder.v(154)
    wire [1:0]\oc8051_top_1/oc8051_decoder1/wr_sfr ;   // oc8051_decoder.v(153)
    wire [3:0]\oc8051_top_1/oc8051_decoder1/alu_op ;   // oc8051_decoder.v(152)
    wire [7:0]\oc8051_top_1/sub_result ;   // oc8051_top.v(468)
    wire \oc8051_top_1/leave_su_mode ;   // oc8051_top.v(424)
    wire \oc8051_top_1/enter_su_mode ;   // oc8051_top.v(423)
    wire [1:0]\oc8051_top_1/decoder_state ;   // oc8051_top.v(258)
    wire [31:0]\oc8051_top_1/idat_i ;   // oc8051_top.v(418)
    wire \oc8051_top_1/istb_o ;   // oc8051_top.v(416)
    wire \oc8051_top_1/iack_i ;   // oc8051_top.v(415)
    wire \oc8051_top_1/bit_addr_o ;   // oc8051_top.v(410)
    wire \oc8051_top_1/bit_out ;   // oc8051_top.v(409)
    wire \oc8051_top_1/bit_data ;   // oc8051_top.v(408)
    wire \oc8051_top_1/bit_addr ;   // oc8051_top.v(407)
    wire [2:0]\oc8051_top_1/op1_cur ;   // oc8051_top.v(405)
    wire \oc8051_top_1/comp_wait ;   // oc8051_top.v(404)
    wire \oc8051_top_1/wr_ind ;   // oc8051_top.v(403)
    wire \oc8051_top_1/rd_ind ;   // oc8051_top.v(402)
    wire \oc8051_top_1/cy ;   // oc8051_top.v(401)
    wire \oc8051_top_1/srcAc ;   // oc8051_top.v(400)
    wire \oc8051_top_1/eq ;   // oc8051_top.v(399)
    wire [1:0]\oc8051_top_1/comp_sel ;   // oc8051_top.v(398)
    wire [15:0]\oc8051_top_1/pc_log_prev ;   // oc8051_top.v(231)
    wire [15:0]\oc8051_top_1/pc_log ;   // oc8051_top.v(230)
    wire \oc8051_top_1/decoder_new_valid_pc ;   // oc8051_top.v(394)
    wire \oc8051_top_1/irom_out_of_rst ;   // oc8051_top.v(391)
    wire [7:0]\oc8051_top_1/op3_n ;   // oc8051_top.v(390)
    wire [7:0]\oc8051_top_1/op2_n ;   // oc8051_top.v(389)
    wire [7:0]\oc8051_top_1/op1_n ;   // oc8051_top.v(388)
    wire [2:0]\oc8051_top_1/pc_wr_sel ;   // oc8051_top.v(386)
    wire \oc8051_top_1/pc_wr ;   // oc8051_top.v(385)
    wire \oc8051_top_1/rd ;   // oc8051_top.v(384)
    wire \oc8051_top_1/wr_o ;   // oc8051_top.v(382)
    wire \oc8051_top_1/wr ;   // oc8051_top.v(381)
    wire \oc8051_top_1/alu_cy ;   // oc8051_top.v(380)
    wire \oc8051_top_1/desOv ;   // oc8051_top.v(379)
    wire \oc8051_top_1/desAc ;   // oc8051_top.v(378)
    wire \oc8051_top_1/desCy ;   // oc8051_top.v(377)
    wire [7:0]\oc8051_top_1/des2 ;   // oc8051_top.v(376)
    wire [7:0]\oc8051_top_1/des1 ;   // oc8051_top.v(375)
    wire [7:0]\oc8051_top_1/des_acc ;   // oc8051_top.v(374)
    wire [7:0]\oc8051_top_1/src3 ;   // oc8051_top.v(373)
    wire [7:0]\oc8051_top_1/src2 ;   // oc8051_top.v(372)
    wire [7:0]\oc8051_top_1/src1 ;   // oc8051_top.v(371)
    wire [1:0]\oc8051_top_1/psw_set ;   // oc8051_top.v(369)
    wire [3:0]\oc8051_top_1/alu_op ;   // oc8051_top.v(368)
    wire [2:0]\oc8051_top_1/mem_act ;   // oc8051_top.v(367)
    wire [7:0]\oc8051_top_1/int_src ;   // oc8051_top.v(364)
    wire \oc8051_top_1/istb ;   // oc8051_top.v(363)
    wire \oc8051_top_1/int_ack ;   // oc8051_top.v(362)
    wire \oc8051_top_1/intr ;   // oc8051_top.v(361)
    wire \oc8051_top_1/reti ;   // oc8051_top.v(360)
    wire \oc8051_top_1/ea_int ;   // oc8051_top.v(358)
    wire \oc8051_top_1/rmw ;   // oc8051_top.v(357)
    wire [1:0]\oc8051_top_1/bank_sel ;   // oc8051_top.v(355)
    wire [1:0]\oc8051_top_1/cy_sel ;   // oc8051_top.v(354)
    wire \oc8051_top_1/sfr_bit ;   // oc8051_top.v(352)
    wire [7:0]\oc8051_top_1/rd_addr ;   // oc8051_top.v(351)
    wire [7:0]\oc8051_top_1/wr_addr ;   // oc8051_top.v(350)
    wire [7:0]\oc8051_top_1/wr_dat ;   // oc8051_top.v(349)
    wire [7:0]\oc8051_top_1/sfr_out ;   // oc8051_top.v(348)
    wire [7:0]\oc8051_top_1/ram_out ;   // oc8051_top.v(347)
    wire [7:0]\oc8051_top_1/ram_data ;   // oc8051_top.v(346)
    wire [2:0]\oc8051_top_1/src_sel1 ;   // oc8051_top.v(344)
    wire [2:0]\oc8051_top_1/ram_wr_sel ;   // oc8051_top.v(343)
    wire [2:0]\oc8051_top_1/ram_rd_sel ;   // oc8051_top.v(342)
    wire [1:0]\oc8051_top_1/src_sel2 ;   // oc8051_top.v(341)
    wire [1:0]\oc8051_top_1/wr_sfr ;   // oc8051_top.v(340)
    wire \oc8051_top_1/src_sel3 ;   // oc8051_top.v(339)
    wire [15:0]\oc8051_top_1/etr ;   // oc8051_top.v(335)
    wire [15:0]\oc8051_top_1/mem_pc ;   // oc8051_top.v(334)
    wire [15:0]\oc8051_top_1/pc ;   // oc8051_top.v(228)
    wire [31:0]\oc8051_top_1/idat_onchip ;   // oc8051_top.v(330)
    wire [7:0]\oc8051_top_1/sp_w ;   // oc8051_top.v(328)
    wire [7:0]\oc8051_top_1/sp ;   // oc8051_top.v(234)
    wire [7:0]\oc8051_top_1/b_reg ;   // oc8051_top.v(236)
    wire [7:0]\oc8051_top_1/acc ;   // oc8051_top.v(235)
    wire [7:0]\oc8051_top_1/op3 ;   // oc8051_top.v(239)
    wire [7:0]\oc8051_top_1/op2 ;   // oc8051_top.v(239)
    wire \oc8051_top_1/oc8051_decoder1/wr ;   // oc8051_decoder.v(151)
    wire [7:0]\oc8051_top_1/op1_d ;   // oc8051_top.v(239)
    wire [7:0]\oc8051_top_1/op1 ;   // oc8051_top.v(239)
    wire [7:0]\oc8051_top_1/ri ;   // oc8051_top.v(316)
    wire [7:0]\oc8051_top_1/dptr_lo ;   // oc8051_top.v(315)
    wire [7:0]\oc8051_top_1/dptr_hi ;   // oc8051_top.v(314)
    wire [15:0]\oc8051_top_1/wbi_adr_o ;   // oc8051_top.v(254)
    wire \oc8051_top_1/wbi_cyc_o ;   // oc8051_top.v(249)
    wire \oc8051_top_1/wbi_stb_o ;   // oc8051_top.v(248)
    wire [7:0]\oc8051_top_1/ie ;   // oc8051_top.v(240)
    wire [2047:0]\oc8051_top_1/iram ;   // oc8051_top.v(238)
    wire [0:1]ea;   // oc8051_tb.v(134)
    wire [15:0]cxrom_addr;   // oc8051_tb.v(142)
    wire [31:0]cxrom_data_out;   // oc8051_tb.v(143)
    wire \oc8051_top_1/p ;   // oc8051_top.v(233)
    wire [7:0]\oc8051_top_1/psw ;   // oc8051_top.v(232)
    wire [2047:0]\oc8051_xiommu1/exp_n ;   // oc8051_xiommu.v(67)
    wire \oc8051_xiommu1/proc_stb ;   // oc8051_xiommu.v(84)
    wire \oc8051_xiommu1/proc_ack ;   // oc8051_xiommu.v(84)
    wire \oc8051_xiommu1/proc_wr ;   // oc8051_xiommu.v(84)
    wire [15:0]\oc8051_xiommu1/proc_addr ;   // oc8051_xiommu.v(86)
    wire [15:0]\oc8051_xiommu1/dpc_ot ;   // oc8051_xiommu.v(86)
    wire [7:0]\oc8051_xiommu1/proc_data_in ;   // oc8051_xiommu.v(87)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbit_winner ;   // oc8051_procarbiter.v(128)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_next ;   // oc8051_procarbiter.v(118)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_inuse_next ;   // oc8051_procarbiter.v(111)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/ack_A ;   // oc8051_procarbiter.v(53)
    wire \oc8051_xiommu1/proc0_ack ;   // oc8051_xiommu.v(60)
    wire [7:0]\oc8051_xiommu1/proc0_data_out ;   // oc8051_xiommu.v(58)
    wire [2:0]\oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next ;   // oc8051_memarbiter.v(185)
    wire [2:0]\oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder ;   // oc8051_memarbiter.v(123)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder_next ;   // oc8051_procarbiter.v(138)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_idle_next ;   // oc8051_procarbiter.v(114)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/ack_B ;   // oc8051_procarbiter.v(63)
    wire \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder ;   // oc8051_procarbiter.v(87)
    wire [7:0]\oc8051_xiommu1/data_out_aes ;   // oc8051_xiommu.v(125)
    wire [7:0]\oc8051_xiommu1/data_out_sha ;   // oc8051_xiommu.v(126)
    wire [7:0]\oc8051_xiommu1/data_out_exp ;   // oc8051_xiommu.v(127)
    wire [7:0]\oc8051_xiommu1/data_out_memwr ;   // oc8051_xiommu.v(128)
    wire [7:0]\oc8051_xiommu1/data_out_pt ;   // oc8051_xiommu.v(129)
    wire [7:0]\oc8051_xiommu1/data_out_ia ;   // oc8051_xiommu.v(130)
    wire [15:0]\oc8051_xiommu1/aes_xram_addr ;   // oc8051_xiommu.v(147)
    wire [7:0]\oc8051_xiommu1/aes_xram_data_out ;   // oc8051_xiommu.v(148)
    wire [7:0]\oc8051_xiommu1/aes_xram_data_in ;   // oc8051_xiommu.v(149)
    wire \oc8051_xiommu1/aes_xram_stb ;   // oc8051_xiommu.v(151)
    wire [15:0]\oc8051_xiommu1/sha_xram_addr ;   // oc8051_xiommu.v(180)
    wire [7:0]\oc8051_xiommu1/sha_xram_data_out ;   // oc8051_xiommu.v(181)
    wire \oc8051_xiommu1/sha_xram_ack ;   // oc8051_xiommu.v(183)
    wire \oc8051_xiommu1/sha_xram_stb ;   // oc8051_xiommu.v(184)
    wire \oc8051_xiommu1/sha_xram_wr ;   // oc8051_xiommu.v(185)
    wire [15:0]\oc8051_xiommu1/exp_xram_addr ;   // oc8051_xiommu.v(212)
    wire [7:0]\oc8051_xiommu1/exp_xram_data_out ;   // oc8051_xiommu.v(213)
    wire \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_next ;   // oc8051_memarbiter.v(170)
    wire \oc8051_xiommu1/exp_xram_ack ;   // oc8051_xiommu.v(215)
    wire \oc8051_xiommu1/exp_xram_stb ;   // oc8051_xiommu.v(216)
    wire \oc8051_xiommu1/exp_xram_wr ;   // oc8051_xiommu.v(217)
    wire [15:0]\oc8051_xiommu1/memwr_xram_addr ;   // oc8051_xiommu.v(244)
    wire [7:0]\oc8051_xiommu1/memwr_xram_data_out ;   // oc8051_xiommu.v(245)
    wire [2:0]\oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner ;   // oc8051_memarbiter.v(179)
    wire \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_idle_next ;   // oc8051_memarbiter.v(167)
    wire \oc8051_xiommu1/memwr_xram_ack ;   // oc8051_xiommu.v(247)
    wire \oc8051_xiommu1/memwr_xram_stb ;   // oc8051_xiommu.v(248)
    wire \oc8051_xiommu1/memwr_xram_wr ;   // oc8051_xiommu.v(249)
    wire \oc8051_xiommu1/stb_out ;   // oc8051_xiommu.v(305)
    wire \oc8051_xiommu1/ack_in ;   // oc8051_xiommu.v(305)
    wire \oc8051_xiommu1/wr_out ;   // oc8051_xiommu.v(305)
    wire [2:0]\oc8051_xiommu1/selected_port ;   // oc8051_xiommu.v(306)
    wire [15:0]\oc8051_xiommu1/addr_out ;   // oc8051_xiommu.v(307)
    wire [7:0]\oc8051_xiommu1/memarbiter_data_in ;   // oc8051_xiommu.v(308)
    wire \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_inuse_next ;   // oc8051_memarbiter.v(164)
    wire \oc8051_xiommu1/aes_top_i/sel_reg_start ;   // aes_top.v(97)
    wire \oc8051_xiommu1/aes_top_i/wren ;   // aes_top.v(126)
    wire \oc8051_xiommu1/aes_top_i/aes_reg_keysel_next ;   // aes_top.v(131)
    wire [7:0]\oc8051_xiommu1/aes_top_i/aes_addr_dataout ;   // aes_top.v(135)
    wire [7:0]\oc8051_xiommu1/aes_top_i/aes_len_dataout ;   // aes_top.v(149)
    wire [7:0]\oc8051_xiommu1/aes_top_i/aes_ctr_dataout ;   // aes_top.v(166)
    wire [7:0]\oc8051_xiommu1/aes_top_i/aes_key0_dataout ;   // aes_top.v(180)
    wire [7:0]\oc8051_xiommu1/aes_top_i/aes_key1_dataout ;   // aes_top.v(194)
    wire [15:0]\oc8051_xiommu1/aes_top_i/operated_bytes_count ;   // aes_top.v(211)
    wire [15:0]\oc8051_xiommu1/aes_top_i/operated_bytes_count_next ;   // aes_top.v(212)
    wire [15:0]\oc8051_xiommu1/aes_top_i/block_counter ;   // aes_top.v(218)
    wire [15:0]\oc8051_xiommu1/aes_top_i/block_counter_next ;   // aes_top.v(219)
    wire [3:0]\oc8051_xiommu1/aes_top_i/byte_counter ;   // aes_top.v(224)
    wire [3:0]\oc8051_xiommu1/aes_top_i/byte_counter_next ;   // aes_top.v(227)
    wire [1:0]\oc8051_xiommu1/aes_top_i/aes_reg_state_next_read_data ;   // aes_top.v(243)
    wire [1:0]\oc8051_xiommu1/aes_top_i/aes_reg_state_next_write_data ;   // aes_top.v(245)
    wire [1:0]\oc8051_xiommu1/aes_top_i/aes_reg_state_next ;   // aes_top.v(251)
    wire [127:0]\oc8051_xiommu1/aes_top_i/mem_data_buf ;   // aes_top.v(261)
    wire [127:0]\oc8051_xiommu1/aes_top_i/mem_data_buf_next ;   // aes_top.v(262)
    wire [127:0]\oc8051_xiommu1/aes_top_i/aes_ctr_v ;   // aes_top.v(281)
    wire [127:0]\oc8051_xiommu1/aes_top_i/aes_out ;   // aes_top.v(282)
    wire [127:0]\oc8051_xiommu1/aes_top_i/encrypted_data ;   // aes_top.v(283)
    wire [127:0]\oc8051_xiommu1/aes_top_i/aes_curr_key ;   // aes_top.v(284)
    wire [127:0]\oc8051_xiommu1/aes_top_i/encrypted_data_buf ;   // aes_top.v(294)
    wire [127:0]\oc8051_xiommu1/aes_top_i/encrypted_data_buf_next ;   // aes_top.v(295)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] ;   // oc8051_page_table.v(44)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] ;   // oc8051_page_table.v(45)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/data_out_wr ;   // oc8051_page_table.v(50)
    wire [7:0]\oc8051_xiommu1/oc8051_page_table_i/data_out_rd ;   // oc8051_page_table.v(50)
    wire [15:0]\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg ;   // oc8051_page_table.v(119)
    wire [1:0]\oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg ;   // oc8051_page_table.v(120)
    wire [2:0]\oc8051_xiommu1/oc8051_page_table_i/illegal_src ;   // oc8051_page_table.v(121)
    wire [15:0]\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg ;   // oc8051_page_table.v(122)
    wire \oc8051_xiommu1/oc8051_page_table_i/accesser ;   // oc8051_page_table.v(129)
    wire [15:0]\oc8051_xiommu1/oc8051_page_table_i/ia_reg_next ;   // oc8051_page_table.v(132)
    wire [2:0]\oc8051_xiommu1/oc8051_page_table_i/ia_src_next ;   // oc8051_page_table.v(133)
    wire \oc8051_xiommu1/oc8051_page_table_i/ia_pc_hi ;   // oc8051_page_table.v(74)
    
    wire \oc8051_top_1/oc8051_decoder1/n1424 , \oc8051_top_1/oc8051_decoder1/n1423 , 
        \oc8051_top_1/oc8051_decoder1/n1422 , \oc8051_top_1/oc8051_decoder1/n1421 , 
        \oc8051_top_1/oc8051_decoder1/n1420 , \oc8051_top_1/oc8051_decoder1/n1419 , 
        \oc8051_top_1/oc8051_decoder1/n1418 , \oc8051_top_1/oc8051_decoder1/n1367 , 
        \oc8051_top_1/oc8051_decoder1/n1366 , \oc8051_top_1/oc8051_decoder1/n1365 , 
        \oc8051_top_1/oc8051_decoder1/n1364 , \oc8051_top_1/oc8051_decoder1/n1363 , 
        \oc8051_top_1/oc8051_decoder1/n1362 , \oc8051_top_1/oc8051_decoder1/n1361 , 
        \oc8051_top_1/oc8051_decoder1/n1360 , \oc8051_top_1/oc8051_decoder1/n1358 , 
        \oc8051_top_1/oc8051_decoder1/n1354 , \oc8051_top_1/oc8051_decoder1/n1351 , 
        \oc8051_top_1/oc8051_decoder1/n1348 , \oc8051_top_1/oc8051_decoder1/n1344 , 
        \oc8051_top_1/oc8051_decoder1/n1341 , \oc8051_top_1/oc8051_decoder1/n1338 , 
        \oc8051_top_1/oc8051_decoder1/n1332 , \oc8051_top_1/oc8051_decoder1/n1330 , 
        \oc8051_top_1/oc8051_decoder1/n1328 , \oc8051_top_1/oc8051_decoder1/n1326 , 
        \oc8051_top_1/oc8051_decoder1/n1324 , \oc8051_top_1/oc8051_decoder1/n1320 , 
        \oc8051_top_1/oc8051_decoder1/n1317 , \oc8051_top_1/oc8051_decoder1/n1312 , 
        \oc8051_top_1/oc8051_decoder1/n1308 , \oc8051_top_1/oc8051_decoder1/n1302 , 
        \oc8051_top_1/oc8051_decoder1/n1297 , \oc8051_top_1/oc8051_decoder1/n1293 , 
        \oc8051_top_1/oc8051_decoder1/n1288 , \oc8051_top_1/oc8051_decoder1/n1283 , 
        \oc8051_top_1/oc8051_decoder1/n1280 , \oc8051_top_1/oc8051_decoder1/n1274 , 
        \oc8051_top_1/oc8051_decoder1/n1272 , \oc8051_top_1/oc8051_decoder1/n1269 , 
        \oc8051_top_1/oc8051_decoder1/n1267 , \oc8051_top_1/oc8051_decoder1/n1262 , 
        \oc8051_top_1/oc8051_decoder1/n1256 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/oc8051_decoder1/n1251 , \oc8051_top_1/oc8051_decoder1/n1250 , 
        \oc8051_top_1/oc8051_decoder1/n1249 , \oc8051_top_1/oc8051_decoder1/n1248 , 
        \oc8051_top_1/oc8051_decoder1/n1246 , \oc8051_top_1/oc8051_decoder1/n1245 , 
        \oc8051_top_1/oc8051_decoder1/n1243 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1241 , \oc8051_top_1/oc8051_decoder1/n1228 , 
        \oc8051_top_1/oc8051_decoder1/n1227 , \oc8051_top_1/oc8051_decoder1/n1226 , 
        \oc8051_top_1/oc8051_decoder1/n1225 , \oc8051_top_1/oc8051_decoder1/n1224 , 
        \oc8051_top_1/oc8051_decoder1/n1223 , \oc8051_top_1/oc8051_decoder1/n1222 , 
        \oc8051_top_1/oc8051_decoder1/n1221 , \oc8051_top_1/oc8051_decoder1/n1198 , 
        \oc8051_top_1/oc8051_decoder1/n1197 , \oc8051_top_1/oc8051_decoder1/n1196 , 
        \oc8051_top_1/oc8051_decoder1/n1195 , \oc8051_top_1/oc8051_decoder1/n1194 , 
        \oc8051_top_1/oc8051_decoder1/n1193 , \oc8051_top_1/oc8051_decoder1/n1192 , 
        \oc8051_top_1/oc8051_decoder1/n1191 , \oc8051_top_1/oc8051_decoder1/n1190 , 
        \oc8051_top_1/oc8051_decoder1/n1189 , \oc8051_top_1/oc8051_decoder1/n1188 , 
        \oc8051_top_1/oc8051_decoder1/n1187 , \oc8051_top_1/oc8051_decoder1/n1186 , 
        \oc8051_top_1/oc8051_decoder1/n1185 , \oc8051_top_1/oc8051_decoder1/n1184 , 
        \oc8051_top_1/oc8051_decoder1/n1183 , \oc8051_top_1/oc8051_decoder1/n1182 , 
        \oc8051_top_1/oc8051_decoder1/n1181 , \oc8051_top_1/oc8051_decoder1/n1180 , 
        \oc8051_top_1/oc8051_decoder1/n1179 , \oc8051_top_1/oc8051_decoder1/n1178 , 
        \oc8051_top_1/oc8051_decoder1/n1177 , \oc8051_top_1/oc8051_decoder1/n1176 , 
        \oc8051_top_1/oc8051_decoder1/n1175 , \oc8051_top_1/oc8051_decoder1/n1174 , 
        \oc8051_top_1/oc8051_decoder1/n1173 , \oc8051_top_1/oc8051_decoder1/n1172 , 
        \oc8051_top_1/oc8051_decoder1/n1171 , \oc8051_top_1/oc8051_decoder1/n1170 , 
        \oc8051_top_1/oc8051_decoder1/n1169 , \oc8051_top_1/oc8051_decoder1/n1168 , 
        \oc8051_top_1/oc8051_decoder1/n1167 , \oc8051_top_1/oc8051_decoder1/n1166 , 
        \oc8051_top_1/oc8051_decoder1/n1165 , \oc8051_top_1/oc8051_decoder1/n1164 , 
        \oc8051_top_1/oc8051_decoder1/n1163 , \oc8051_top_1/oc8051_decoder1/n1162 , 
        \oc8051_top_1/oc8051_decoder1/n1161 , \oc8051_top_1/oc8051_decoder1/n1160 , 
        \oc8051_top_1/oc8051_decoder1/n1159 , \oc8051_top_1/oc8051_decoder1/n1158 , 
        \oc8051_top_1/oc8051_decoder1/n1157 , \oc8051_top_1/oc8051_decoder1/n1156 , 
        \oc8051_top_1/oc8051_decoder1/n1155 , \oc8051_top_1/oc8051_decoder1/n1154 , 
        \oc8051_top_1/oc8051_decoder1/n1153 , \oc8051_top_1/oc8051_decoder1/n1152 , 
        \oc8051_top_1/oc8051_decoder1/n1151 , \oc8051_top_1/oc8051_decoder1/n1150 , 
        \oc8051_top_1/oc8051_decoder1/n1149 , \oc8051_top_1/oc8051_decoder1/n1148 , 
        \oc8051_top_1/oc8051_decoder1/n1147 , \oc8051_top_1/oc8051_decoder1/n1146 , 
        \oc8051_top_1/oc8051_decoder1/n1145 , \oc8051_top_1/oc8051_decoder1/n1144 , 
        \oc8051_top_1/oc8051_decoder1/n1143 , \oc8051_top_1/oc8051_decoder1/n1142 , 
        \oc8051_top_1/oc8051_decoder1/n1141 , \oc8051_top_1/oc8051_decoder1/n1140 , 
        \oc8051_top_1/oc8051_decoder1/n1129 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1115 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1107 , \oc8051_top_1/oc8051_decoder1/n1095 , 
        \oc8051_top_1/oc8051_decoder1/n1089 , \oc8051_top_1/oc8051_decoder1/n1085 , 
        \oc8051_top_1/oc8051_decoder1/n1082 , \oc8051_top_1/oc8051_decoder1/n1077 , 
        \oc8051_top_1/oc8051_decoder1/n1044 , \oc8051_top_1/oc8051_decoder1/n1015 , 
        \oc8051_top_1/oc8051_decoder1/n1004 , \oc8051_top_1/oc8051_decoder1/n994 , 
        \oc8051_top_1/oc8051_decoder1/n987 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n936 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n922 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/n915 , \oc8051_top_1/oc8051_decoder1/n905 , 
        \oc8051_top_1/oc8051_decoder1/n899 , \oc8051_top_1/oc8051_decoder1/n889 , 
        \oc8051_top_1/oc8051_decoder1/n884 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 , \oc8051_top_1/oc8051_decoder1/n852 , 
        \oc8051_top_1/oc8051_decoder1/n848 , \oc8051_top_1/oc8051_decoder1/n843 , 
        \oc8051_top_1/oc8051_decoder1/n839 , \oc8051_top_1/oc8051_decoder1/n834 , 
        \oc8051_top_1/oc8051_decoder1/n831 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n791 , \oc8051_top_1/oc8051_decoder1/n780 , 
        \oc8051_top_1/oc8051_decoder1/n763 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n750 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n740 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n728 , \oc8051_top_1/oc8051_decoder1/n718 , 
        \oc8051_top_1/oc8051_decoder1/n709 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/n691 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/n679 , \oc8051_top_1/oc8051_decoder1/n675 , 
        \oc8051_top_1/oc8051_decoder1/n643 , \oc8051_top_1/oc8051_decoder1/n642 , 
        \oc8051_top_1/oc8051_decoder1/n641 , \oc8051_top_1/oc8051_decoder1/n640 , 
        \oc8051_top_1/oc8051_decoder1/n613 , \oc8051_top_1/oc8051_decoder1/n612 , 
        \oc8051_top_1/oc8051_decoder1/n611 , \oc8051_top_1/oc8051_decoder1/n607 , 
        \oc8051_top_1/oc8051_decoder1/n565 , \oc8051_top_1/oc8051_decoder1/n564 , 
        \oc8051_top_1/oc8051_decoder1/n563 , \oc8051_top_1/oc8051_decoder1/n561 , 
        \oc8051_top_1/oc8051_decoder1/n560 , \oc8051_top_1/oc8051_decoder1/n559 , 
        \oc8051_top_1/oc8051_decoder1/n558 , \oc8051_top_1/oc8051_decoder1/n557 , 
        \oc8051_top_1/oc8051_decoder1/n556 , \oc8051_top_1/oc8051_decoder1/n555 , 
        \oc8051_top_1/oc8051_decoder1/n553 , \oc8051_top_1/oc8051_decoder1/n552 , 
        \oc8051_top_1/oc8051_decoder1/n551 , \oc8051_top_1/oc8051_decoder1/n550 , 
        \oc8051_top_1/oc8051_decoder1/n549 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n543 , \oc8051_top_1/oc8051_decoder1/n539 , 
        \oc8051_top_1/oc8051_decoder1/n524 , \oc8051_top_1/oc8051_decoder1/n512 , 
        \oc8051_top_1/oc8051_decoder1/n509 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/n502 , \oc8051_top_1/oc8051_decoder1/n497 , 
        \oc8051_top_1/oc8051_decoder1/n493 , \oc8051_top_1/oc8051_decoder1/n490 , 
        \oc8051_top_1/oc8051_decoder1/n482 , \oc8051_top_1/oc8051_decoder1/n477 , 
        \oc8051_top_1/oc8051_decoder1/n473 , \oc8051_top_1/oc8051_decoder1/n469 , 
        \oc8051_top_1/oc8051_decoder1/n464 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n456 , \oc8051_top_1/oc8051_decoder1/n452 , 
        \oc8051_top_1/oc8051_decoder1/n446 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/n436 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n425 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/n402 , \oc8051_top_1/oc8051_decoder1/n397 , 
        \oc8051_top_1/oc8051_decoder1/n382 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n348 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/n323 , \oc8051_top_1/oc8051_decoder1/n317 , 
        \oc8051_top_1/oc8051_decoder1/n312 , \oc8051_top_1/oc8051_decoder1/n307 , 
        \oc8051_top_1/oc8051_decoder1/n303 , \oc8051_top_1/oc8051_decoder1/n270 , 
        \oc8051_top_1/oc8051_decoder1/n258 , \oc8051_top_1/oc8051_decoder1/n255 , 
        \oc8051_top_1/oc8051_decoder1/n252 , \oc8051_top_1/oc8051_decoder1/n248 , 
        \oc8051_top_1/oc8051_decoder1/n241 , \oc8051_top_1/oc8051_decoder1/n217 , 
        \oc8051_top_1/oc8051_decoder1/n215 , \oc8051_top_1/oc8051_decoder1/n209 , 
        \oc8051_top_1/oc8051_decoder1/n208 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/n159 , \oc8051_top_1/oc8051_decoder1/n158 , 
        \oc8051_top_1/oc8051_decoder1/n157 , \oc8051_top_1/oc8051_decoder1/n156 , 
        \oc8051_top_1/oc8051_decoder1/n155 , \oc8051_top_1/oc8051_decoder1/n154 , 
        \oc8051_top_1/oc8051_decoder1/n153 , \oc8051_top_1/oc8051_decoder1/n152 , 
        \oc8051_top_1/oc8051_decoder1/n151 , \oc8051_top_1/oc8051_decoder1/n150 , 
        \oc8051_top_1/oc8051_decoder1/n149 , \oc8051_top_1/oc8051_decoder1/n148 , 
        \oc8051_top_1/oc8051_decoder1/n147 , \oc8051_top_1/oc8051_decoder1/n146 , 
        \oc8051_top_1/oc8051_decoder1/n145 , \oc8051_top_1/oc8051_decoder1/n144 , 
        \oc8051_top_1/oc8051_decoder1/n143 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n127 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n101 , \oc8051_top_1/oc8051_decoder1/n95 , 
        \oc8051_top_1/oc8051_decoder1/n91 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/n84 , \oc8051_top_1/oc8051_decoder1/n83 , 
        \oc8051_top_1/oc8051_decoder1/n80 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/n74 , \oc8051_top_1/oc8051_decoder1/n73 , 
        \oc8051_top_1/oc8051_decoder1/n72 , \oc8051_top_1/oc8051_decoder1/n71 , 
        \oc8051_top_1/oc8051_decoder1/n61 , \oc8051_top_1/oc8051_decoder1/n60 , 
        \oc8051_top_1/oc8051_decoder1/n59 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/n53 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/oc8051_decoder1/n37 , \oc8051_top_1/oc8051_decoder1/n36 , 
        \oc8051_top_1/oc8051_decoder1/n32 , \oc8051_top_1/oc8051_decoder1/n23 , 
        \oc8051_top_1/oc8051_decoder1/n22 , \oc8051_top_1/oc8051_decoder1/n21 , 
        \oc8051_top_1/oc8051_decoder1/n20 , \oc8051_top_1/oc8051_decoder1/n19 , 
        \oc8051_top_1/oc8051_decoder1/n18 , \oc8051_top_1/oc8051_decoder1/n17 , 
        \oc8051_top_1/oc8051_decoder1/n16 , \oc8051_top_1/oc8051_decoder1/n14 , 
        \oc8051_top_1/oc8051_decoder1/n13 , \oc8051_top_1/oc8051_decoder1/n6 , 
        \oc8051_top_1/oc8051_decoder1/n5 , \oc8051_top_1/oc8051_decoder1/n4 , 
        \oc8051_top_1/n78 , \oc8051_top_1/n77 , \oc8051_top_1/n76 , \oc8051_top_1/n72 , 
        \oc8051_top_1/n71 , \oc8051_top_1/n70 , n153, \oc8051_xiommu1/oc8051_procarbiter_i/n67 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n58 , \oc8051_xiommu1/oc8051_memarbiter_i/n43 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n38 , \oc8051_xiommu1/oc8051_memarbiter_i/n14 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n69 , \oc8051_xiommu1/oc8051_procarbiter_i/n64 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n47 , \oc8051_xiommu1/oc8051_memarbiter_i/n42 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n37 , \oc8051_xiommu1/oc8051_memarbiter_i/n13 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n46 , \oc8051_xiommu1/oc8051_memarbiter_i/n41 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n36 , \oc8051_xiommu1/oc8051_memarbiter_i/n26 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n12 , \oc8051_xiommu1/oc8051_memarbiter_i/n45 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n40 , \oc8051_xiommu1/oc8051_memarbiter_i/n25 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n7 , \oc8051_xiommu1/oc8051_memarbiter_i/n44 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n39 , \oc8051_xiommu1/oc8051_memarbiter_i/n24 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n5 , \oc8051_xiommu1/n10 , \oc8051_xiommu1/n11 , 
        \oc8051_xiommu1/n12 , \oc8051_xiommu1/n13 , \oc8051_xiommu1/n14 , 
        \oc8051_xiommu1/n15 , \oc8051_xiommu1/n31 , \oc8051_xiommu1/n32 , 
        \oc8051_xiommu1/n33 , \oc8051_xiommu1/n34 , \oc8051_xiommu1/n35 , 
        \oc8051_xiommu1/n36 , \oc8051_xiommu1/n45 , \oc8051_xiommu1/n47 , 
        \oc8051_xiommu1/n48 , \oc8051_xiommu1/n49 , \oc8051_xiommu1/n50 , 
        \oc8051_xiommu1/n51 , \oc8051_xiommu1/n52 , \oc8051_xiommu1/n53 , 
        \oc8051_xiommu1/n54 , \oc8051_xiommu1/n55 , \oc8051_xiommu1/n56 , 
        \oc8051_xiommu1/n57 , \oc8051_xiommu1/n58 , \oc8051_xiommu1/n59 , 
        \oc8051_xiommu1/n60 , \oc8051_xiommu1/n61 , \oc8051_xiommu1/n62 , 
        \oc8051_xiommu1/n63 , \oc8051_xiommu1/n64 , \oc8051_xiommu1/n65 , 
        \oc8051_xiommu1/n66 , \oc8051_xiommu1/n67 , \oc8051_xiommu1/n68 , 
        \oc8051_xiommu1/n69 , \oc8051_xiommu1/n70 , \oc8051_xiommu1/n71 , 
        \oc8051_xiommu1/n72 , \oc8051_xiommu1/n73 , \oc8051_xiommu1/n74 , 
        \oc8051_xiommu1/n75 , \oc8051_xiommu1/n76 , \oc8051_xiommu1/n77 , 
        \oc8051_xiommu1/n78 , \oc8051_xiommu1/n79 , \oc8051_xiommu1/n80 , 
        \oc8051_xiommu1/n81 , \oc8051_xiommu1/n82 , \oc8051_xiommu1/n83 , 
        \oc8051_xiommu1/n84 , \oc8051_xiommu1/n85 , \oc8051_xiommu1/n86 , 
        \oc8051_xiommu1/n95 , \oc8051_xiommu1/n96 , \oc8051_xiommu1/n97 , 
        \oc8051_xiommu1/n98 , \oc8051_xiommu1/n99 , \oc8051_xiommu1/n100 , 
        \oc8051_xiommu1/n101 , \oc8051_xiommu1/n102 , \oc8051_xiommu1/n103 , 
        \oc8051_xiommu1/n104 , \oc8051_xiommu1/n105 , \oc8051_xiommu1/n106 , 
        \oc8051_xiommu1/n107 , \oc8051_xiommu1/n108 , \oc8051_xiommu1/n109 , 
        \oc8051_xiommu1/n110 , \oc8051_xiommu1/n111 , \oc8051_xiommu1/n112 , 
        \oc8051_xiommu1/n113 , \oc8051_xiommu1/n114 , \oc8051_xiommu1/n115 , 
        \oc8051_xiommu1/n116 , \oc8051_xiommu1/n117 , \oc8051_xiommu1/n118 , 
        \oc8051_xiommu1/n119 , \oc8051_xiommu1/n120 , \oc8051_xiommu1/n121 , 
        \oc8051_xiommu1/n122 , \oc8051_xiommu1/n123 , \oc8051_xiommu1/n124 , 
        \oc8051_xiommu1/n125 , \oc8051_xiommu1/n126 , \oc8051_xiommu1/n127 , 
        \oc8051_xiommu1/n128 , \oc8051_xiommu1/n129 , \oc8051_xiommu1/n130 , 
        \oc8051_xiommu1/n131 , \oc8051_xiommu1/n132 , \oc8051_xiommu1/n133 , 
        \oc8051_xiommu1/n134 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_58/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n9 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n11 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n13 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n15 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n17 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_144/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_144/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_144/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_144/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_145/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_145/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_145/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_145/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_147/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_147/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_148/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_148/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_150/n1 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n1 , \oc8051_top_1/oc8051_decoder1/Select_151/n2 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n3 , \oc8051_top_1/oc8051_decoder1/Select_151/n4 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n5 , \oc8051_top_1/oc8051_decoder1/Select_151/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_152/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_152/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_152/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_155/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_155/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_155/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_156/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_156/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n8 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n10 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n12 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n14 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n16 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n18 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n20 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n22 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n24 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n26 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n28 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n30 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n32 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n33 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n34 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n35 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n36 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n37 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n38 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n39 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n40 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n41 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n42 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n43 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n44 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n45 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n46 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n47 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n48 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n49 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n50 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n51 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n52 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n53 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n54 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n55 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n56 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n57 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n58 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n59 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n60 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n61 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n62 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n63 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n64 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n65 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n66 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n67 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n68 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n69 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n70 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n71 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n72 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n73 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n74 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n75 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n76 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n77 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n78 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n79 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_549/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_549/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_549/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n28 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n32 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n33 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n35 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_552/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_552/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_552/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n34 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n37 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n38 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n39 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n40 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n41 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n42 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n43 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n44 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n45 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n46 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n47 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n48 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n49 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n50 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n51 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n52 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n53 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n54 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n55 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n57 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n58 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n59 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n60 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n61 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n62 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n63 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n64 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n65 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n66 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n67 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n68 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n69 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n70 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n71 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n72 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n73 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n74 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n75 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n76 , 
        \oc8051_top_1/oc8051_decoder1/Select_556/n1 , \oc8051_top_1/oc8051_decoder1/Select_556/n2 , 
        \oc8051_top_1/oc8051_decoder1/Select_556/n3 , \oc8051_top_1/oc8051_decoder1/Select_556/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_557/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_557/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_557/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_558/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n10 , 
        \oc8051_top_1/oc8051_decoder1/Mux_565/n1 , \oc8051_top_1/oc8051_decoder1/Mux_565/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_566/n1 , \oc8051_top_1/oc8051_decoder1/Mux_566/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_567/n1 , \oc8051_top_1/oc8051_decoder1/Mux_567/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_568/n1 , \oc8051_top_1/oc8051_decoder1/Mux_568/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_569/n1 , \oc8051_top_1/oc8051_decoder1/Mux_569/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_570/n1 , \oc8051_top_1/oc8051_decoder1/Mux_570/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_571/n1 , \oc8051_top_1/oc8051_decoder1/Mux_571/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_572/n1 , \oc8051_top_1/oc8051_decoder1/Mux_572/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_573/n1 , \oc8051_top_1/oc8051_decoder1/Mux_573/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_574/n1 , \oc8051_top_1/oc8051_decoder1/Mux_574/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_575/n1 , \oc8051_top_1/oc8051_decoder1/Mux_575/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_576/n1 , \oc8051_top_1/oc8051_decoder1/Mux_576/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_577/n1 , \oc8051_top_1/oc8051_decoder1/Mux_577/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_578/n1 , \oc8051_top_1/oc8051_decoder1/Mux_578/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_610/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_640/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_641/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1141/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1141/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n34 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n34 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n37 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n38 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n39 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n40 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n41 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n42 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n43 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n28 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n32 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n34 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n28 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n32 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n33 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n35 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n2 , \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n34 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n37 , \oc8051_top_1/oc8051_decoder1/Mux_1158/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1158/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1159/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1159/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1160/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1160/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1161/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1161/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1162/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1162/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1163/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1163/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1164/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1164/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1165/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1165/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1166/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1166/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1167/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1167/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1168/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1168/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1169/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1169/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1170/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1170/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1171/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1171/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1172/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1172/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1173/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1173/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1174/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1174/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1175/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1175/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1176/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1176/n2 , \oc8051_top_1/oc8051_decoder1/Mux_1177/n1 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1177/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1219/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n2 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n8 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n10 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n12 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n14 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n16 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n18 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n20 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n22 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n24 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n26 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n28 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n4 , 
        \oc8051_top_1/oc8051_decoder1/Select_1362/n1 , \oc8051_top_1/oc8051_decoder1/Select_1362/n2 , 
        \oc8051_top_1/oc8051_decoder1/Select_1362/n3 , \oc8051_top_1/oc8051_decoder1/Select_1362/n4 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1363/n1 , \oc8051_top_1/oc8051_decoder1/Mux_1363/n2 , 
        \oc8051_top_1/oc8051_decoder1/Mux_1364/n1 , \oc8051_top_1/oc8051_decoder1/Mux_1364/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n1 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1418/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1419/n1 , \oc8051_top_1/oc8051_decoder1/reduce_or_1420/n1 , 
        \oc8051_xiommu1/aes_top_i/n4 , \oc8051_xiommu1/aes_top_i/n5 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 , \oc8051_xiommu1/aes_top_i/n10 , \oc8051_xiommu1/aes_top_i/n11 , 
        \oc8051_xiommu1/aes_top_i/n12 , \oc8051_xiommu1/aes_top_i/n13 , 
        \oc8051_xiommu1/aes_top_i/n14 , \oc8051_xiommu1/aes_top_i/n15 , 
        \oc8051_xiommu1/aes_top_i/n17 , \oc8051_xiommu1/aes_top_i/n27 , 
        \oc8051_xiommu1/aes_top_i/n28 , \oc8051_xiommu1/aes_top_i/n58 , 
        \oc8051_xiommu1/aes_top_i/n68 , \oc8051_xiommu1/aes_top_i/n89 , 
        \oc8051_xiommu1/aes_top_i/n90 , \oc8051_xiommu1/aes_top_i/n91 , 
        \oc8051_xiommu1/aes_top_i/n92 , \oc8051_xiommu1/aes_top_i/n93 , 
        \oc8051_xiommu1/aes_top_i/n94 , \oc8051_xiommu1/aes_top_i/n95 , 
        \oc8051_xiommu1/aes_top_i/n96 , \oc8051_xiommu1/aes_top_i/n97 , 
        \oc8051_xiommu1/aes_top_i/n98 , \oc8051_xiommu1/aes_top_i/n99 , 
        \oc8051_xiommu1/aes_top_i/n100 , \oc8051_xiommu1/aes_top_i/n101 , 
        \oc8051_xiommu1/aes_top_i/n102 , \oc8051_xiommu1/aes_top_i/n103 , 
        \oc8051_xiommu1/aes_top_i/n104 , \oc8051_xiommu1/aes_top_i/n105 , 
        \oc8051_xiommu1/aes_top_i/n106 , \oc8051_xiommu1/aes_top_i/n107 , 
        \oc8051_xiommu1/aes_top_i/n108 , \oc8051_xiommu1/aes_top_i/n109 , 
        \oc8051_xiommu1/aes_top_i/n110 , \oc8051_xiommu1/aes_top_i/n111 , 
        \oc8051_xiommu1/aes_top_i/n112 , \oc8051_xiommu1/aes_top_i/n113 , 
        \oc8051_xiommu1/aes_top_i/n114 , \oc8051_xiommu1/aes_top_i/n115 , 
        \oc8051_xiommu1/aes_top_i/n116 , \oc8051_xiommu1/aes_top_i/n117 , 
        \oc8051_xiommu1/aes_top_i/n118 , \oc8051_xiommu1/aes_top_i/n119 , 
        \oc8051_xiommu1/aes_top_i/n120 , \oc8051_xiommu1/aes_top_i/n121 , 
        \oc8051_xiommu1/aes_top_i/n122 , \oc8051_xiommu1/aes_top_i/n123 , 
        \oc8051_xiommu1/aes_top_i/n124 , \oc8051_xiommu1/aes_top_i/n125 , 
        \oc8051_xiommu1/aes_top_i/n126 , \oc8051_xiommu1/aes_top_i/n127 , 
        \oc8051_xiommu1/aes_top_i/n128 , \oc8051_xiommu1/aes_top_i/n129 , 
        \oc8051_xiommu1/aes_top_i/n130 , \oc8051_xiommu1/aes_top_i/n131 , 
        \oc8051_xiommu1/aes_top_i/n132 , \oc8051_xiommu1/aes_top_i/n133 , 
        \oc8051_xiommu1/aes_top_i/n134 , \oc8051_xiommu1/aes_top_i/n135 , 
        \oc8051_xiommu1/aes_top_i/n136 , \oc8051_xiommu1/aes_top_i/n146 , 
        \oc8051_xiommu1/aes_top_i/n148 , \oc8051_xiommu1/aes_top_i/n154 , 
        \oc8051_xiommu1/aes_top_i/n158 , \oc8051_xiommu1/aes_top_i/n159 , 
        \oc8051_xiommu1/aes_top_i/n160 , \oc8051_xiommu1/aes_top_i/n161 , 
        \oc8051_xiommu1/aes_top_i/n162 , \oc8051_xiommu1/aes_top_i/n165 , 
        \oc8051_xiommu1/aes_top_i/n166 , \oc8051_xiommu1/aes_top_i/n167 , 
        \oc8051_xiommu1/aes_top_i/n168 , \oc8051_xiommu1/aes_top_i/n169 , 
        \oc8051_xiommu1/aes_top_i/n170 , \oc8051_xiommu1/aes_top_i/n171 , 
        \oc8051_xiommu1/aes_top_i/n172 , \oc8051_xiommu1/aes_top_i/n173 , 
        \oc8051_xiommu1/aes_top_i/n174 , \oc8051_xiommu1/aes_top_i/n175 , 
        \oc8051_xiommu1/aes_top_i/n176 , \oc8051_xiommu1/aes_top_i/n178 , 
        \oc8051_xiommu1/aes_top_i/n179 , \oc8051_xiommu1/aes_top_i/n180 , 
        \oc8051_xiommu1/aes_top_i/n181 , \oc8051_xiommu1/aes_top_i/n182 , 
        \oc8051_xiommu1/aes_top_i/n183 , \oc8051_xiommu1/aes_top_i/n184 , 
        \oc8051_xiommu1/aes_top_i/n185 , \oc8051_xiommu1/aes_top_i/n186 , 
        \oc8051_xiommu1/aes_top_i/n187 , \oc8051_xiommu1/aes_top_i/n188 , 
        \oc8051_xiommu1/aes_top_i/n189 , \oc8051_xiommu1/aes_top_i/n208 , 
        \oc8051_xiommu1/aes_top_i/n209 , \oc8051_xiommu1/aes_top_i/n210 , 
        \oc8051_xiommu1/aes_top_i/n211 , \oc8051_xiommu1/aes_top_i/n212 , 
        \oc8051_xiommu1/aes_top_i/n213 , \oc8051_xiommu1/aes_top_i/n214 , 
        \oc8051_xiommu1/aes_top_i/n215 , \oc8051_xiommu1/aes_top_i/n216 , 
        \oc8051_xiommu1/aes_top_i/n217 , \oc8051_xiommu1/aes_top_i/n218 , 
        \oc8051_xiommu1/aes_top_i/n219 , \oc8051_xiommu1/aes_top_i/n221 , 
        \oc8051_xiommu1/aes_top_i/n222 , \oc8051_xiommu1/aes_top_i/n223 , 
        \oc8051_xiommu1/aes_top_i/n224 , \oc8051_xiommu1/aes_top_i/n225 , 
        \oc8051_xiommu1/aes_top_i/n226 , \oc8051_xiommu1/aes_top_i/n227 , 
        \oc8051_xiommu1/aes_top_i/n228 , \oc8051_xiommu1/aes_top_i/n229 , 
        \oc8051_xiommu1/aes_top_i/n230 , \oc8051_xiommu1/aes_top_i/n231 , 
        \oc8051_xiommu1/aes_top_i/n232 , \oc8051_xiommu1/aes_top_i/n251 , 
        \oc8051_xiommu1/aes_top_i/n252 , \oc8051_xiommu1/aes_top_i/n253 , 
        \oc8051_xiommu1/aes_top_i/n254 , \oc8051_xiommu1/aes_top_i/n256 , 
        \oc8051_xiommu1/aes_top_i/n257 , \oc8051_xiommu1/aes_top_i/n258 , 
        \oc8051_xiommu1/aes_top_i/n259 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/n266 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/n268 , \oc8051_xiommu1/aes_top_i/n269 , 
        \oc8051_xiommu1/aes_top_i/n272 , \oc8051_xiommu1/aes_top_i/n275 , 
        \oc8051_xiommu1/aes_top_i/n276 , \oc8051_xiommu1/aes_top_i/n277 , 
        \oc8051_xiommu1/aes_top_i/n278 , \oc8051_xiommu1/aes_top_i/n279 , 
        \oc8051_xiommu1/aes_top_i/n280 , \oc8051_xiommu1/aes_top_i/n281 , 
        \oc8051_xiommu1/aes_top_i/n282 , \oc8051_xiommu1/aes_top_i/n283 , 
        \oc8051_xiommu1/aes_top_i/n284 , \oc8051_xiommu1/aes_top_i/n285 , 
        \oc8051_xiommu1/aes_top_i/n286 , \oc8051_xiommu1/aes_top_i/n287 , 
        \oc8051_xiommu1/aes_top_i/n288 , \oc8051_xiommu1/aes_top_i/n289 , 
        \oc8051_xiommu1/aes_top_i/n290 , \oc8051_xiommu1/aes_top_i/n315 , 
        \oc8051_xiommu1/aes_top_i/n316 , \oc8051_xiommu1/aes_top_i/n317 , 
        \oc8051_xiommu1/aes_top_i/n318 , \oc8051_xiommu1/aes_top_i/n319 , 
        \oc8051_xiommu1/aes_top_i/n320 , \oc8051_xiommu1/aes_top_i/n323 , 
        \oc8051_xiommu1/aes_top_i/n324 , \oc8051_xiommu1/aes_top_i/n1074 , 
        \oc8051_xiommu1/aes_top_i/n1075 , \oc8051_xiommu1/aes_top_i/n1076 , 
        \oc8051_xiommu1/aes_top_i/n1077 , \oc8051_xiommu1/aes_top_i/n1078 , 
        \oc8051_xiommu1/aes_top_i/n1079 , \oc8051_xiommu1/aes_top_i/n1080 , 
        \oc8051_xiommu1/aes_top_i/n1081 , \oc8051_xiommu1/aes_top_i/n1082 , 
        \oc8051_xiommu1/aes_top_i/n1083 , \oc8051_xiommu1/aes_top_i/n1084 , 
        \oc8051_xiommu1/aes_top_i/n1085 , \oc8051_xiommu1/aes_top_i/n1086 , 
        \oc8051_xiommu1/aes_top_i/n1087 , \oc8051_xiommu1/aes_top_i/n1088 , 
        \oc8051_xiommu1/aes_top_i/n1089 , \oc8051_xiommu1/aes_top_i/n1090 , 
        \oc8051_xiommu1/aes_top_i/n1091 , \oc8051_xiommu1/aes_top_i/n1092 , 
        \oc8051_xiommu1/aes_top_i/n1093 , \oc8051_xiommu1/aes_top_i/n1094 , 
        \oc8051_xiommu1/aes_top_i/n1095 , \oc8051_xiommu1/aes_top_i/n1096 , 
        \oc8051_xiommu1/aes_top_i/n1097 , \oc8051_xiommu1/aes_top_i/n1098 , 
        \oc8051_xiommu1/aes_top_i/n1099 , \oc8051_xiommu1/aes_top_i/n1100 , 
        \oc8051_xiommu1/aes_top_i/n1101 , \oc8051_xiommu1/aes_top_i/n1102 , 
        \oc8051_xiommu1/aes_top_i/n1103 , \oc8051_xiommu1/aes_top_i/n1104 , 
        \oc8051_xiommu1/aes_top_i/n1105 , \oc8051_xiommu1/aes_top_i/n1106 , 
        \oc8051_xiommu1/aes_top_i/n1107 , \oc8051_xiommu1/aes_top_i/n1108 , 
        \oc8051_xiommu1/aes_top_i/n1109 , \oc8051_xiommu1/aes_top_i/n1110 , 
        \oc8051_xiommu1/aes_top_i/n1111 , \oc8051_xiommu1/aes_top_i/n1112 , 
        \oc8051_xiommu1/aes_top_i/n1113 , \oc8051_xiommu1/aes_top_i/n1114 , 
        \oc8051_xiommu1/aes_top_i/n1115 , \oc8051_xiommu1/aes_top_i/n1116 , 
        \oc8051_xiommu1/aes_top_i/n1117 , \oc8051_xiommu1/aes_top_i/n1118 , 
        \oc8051_xiommu1/aes_top_i/n1119 , \oc8051_xiommu1/aes_top_i/n1120 , 
        \oc8051_xiommu1/aes_top_i/n1121 , \oc8051_xiommu1/aes_top_i/n1122 , 
        \oc8051_xiommu1/aes_top_i/n1123 , \oc8051_xiommu1/aes_top_i/n1124 , 
        \oc8051_xiommu1/aes_top_i/n1125 , \oc8051_xiommu1/aes_top_i/n1126 , 
        \oc8051_xiommu1/aes_top_i/n1127 , \oc8051_xiommu1/aes_top_i/n1128 , 
        \oc8051_xiommu1/aes_top_i/n1129 , \oc8051_xiommu1/aes_top_i/n1130 , 
        \oc8051_xiommu1/aes_top_i/n1131 , \oc8051_xiommu1/aes_top_i/n1132 , 
        \oc8051_xiommu1/aes_top_i/n1133 , \oc8051_xiommu1/aes_top_i/n1134 , 
        \oc8051_xiommu1/aes_top_i/n1135 , \oc8051_xiommu1/aes_top_i/n1136 , 
        \oc8051_xiommu1/aes_top_i/n1137 , \oc8051_xiommu1/aes_top_i/n1138 , 
        \oc8051_xiommu1/aes_top_i/n1139 , \oc8051_xiommu1/aes_top_i/n1140 , 
        \oc8051_xiommu1/aes_top_i/n1141 , \oc8051_xiommu1/aes_top_i/n1142 , 
        \oc8051_xiommu1/aes_top_i/n1143 , \oc8051_xiommu1/aes_top_i/n1144 , 
        \oc8051_xiommu1/aes_top_i/n1145 , \oc8051_xiommu1/aes_top_i/n1146 , 
        \oc8051_xiommu1/aes_top_i/n1147 , \oc8051_xiommu1/aes_top_i/n1148 , 
        \oc8051_xiommu1/aes_top_i/n1149 , \oc8051_xiommu1/aes_top_i/n1150 , 
        \oc8051_xiommu1/aes_top_i/n1151 , \oc8051_xiommu1/aes_top_i/n1152 , 
        \oc8051_xiommu1/aes_top_i/n1153 , \oc8051_xiommu1/aes_top_i/n1154 , 
        \oc8051_xiommu1/aes_top_i/n1155 , \oc8051_xiommu1/aes_top_i/n1156 , 
        \oc8051_xiommu1/aes_top_i/n1157 , \oc8051_xiommu1/aes_top_i/n1158 , 
        \oc8051_xiommu1/aes_top_i/n1159 , \oc8051_xiommu1/aes_top_i/n1160 , 
        \oc8051_xiommu1/aes_top_i/n1161 , \oc8051_xiommu1/aes_top_i/n1162 , 
        \oc8051_xiommu1/aes_top_i/n1163 , \oc8051_xiommu1/aes_top_i/n1164 , 
        \oc8051_xiommu1/aes_top_i/n1165 , \oc8051_xiommu1/aes_top_i/n1166 , 
        \oc8051_xiommu1/aes_top_i/n1167 , \oc8051_xiommu1/aes_top_i/n1168 , 
        \oc8051_xiommu1/aes_top_i/n1169 , \oc8051_xiommu1/aes_top_i/n1170 , 
        \oc8051_xiommu1/aes_top_i/n1171 , \oc8051_xiommu1/aes_top_i/n1172 , 
        \oc8051_xiommu1/aes_top_i/n1173 , \oc8051_xiommu1/aes_top_i/n1174 , 
        \oc8051_xiommu1/aes_top_i/n1175 , \oc8051_xiommu1/aes_top_i/n1176 , 
        \oc8051_xiommu1/aes_top_i/n1177 , \oc8051_xiommu1/aes_top_i/n1178 , 
        \oc8051_xiommu1/aes_top_i/n1179 , \oc8051_xiommu1/aes_top_i/n1180 , 
        \oc8051_xiommu1/aes_top_i/n1181 , \oc8051_xiommu1/aes_top_i/n1182 , 
        \oc8051_xiommu1/aes_top_i/n1183 , \oc8051_xiommu1/aes_top_i/n1184 , 
        \oc8051_xiommu1/aes_top_i/n1185 , \oc8051_xiommu1/aes_top_i/n1195 , 
        \oc8051_xiommu1/aes_top_i/n1196 , \oc8051_xiommu1/aes_top_i/n1197 , 
        \oc8051_xiommu1/aes_top_i/n1198 , \oc8051_xiommu1/aes_top_i/n1199 , 
        \oc8051_xiommu1/aes_top_i/n1200 , \oc8051_xiommu1/aes_top_i/n1201 , 
        \oc8051_xiommu1/aes_top_i/n1202 , \oc8051_xiommu1/aes_top_i/n1203 , 
        \oc8051_xiommu1/aes_top_i/n1204 , \oc8051_xiommu1/aes_top_i/n1205 , 
        \oc8051_xiommu1/aes_top_i/n1206 , \oc8051_xiommu1/aes_top_i/n1207 , 
        \oc8051_xiommu1/aes_top_i/n1208 , \oc8051_xiommu1/aes_top_i/n1209 , 
        \oc8051_xiommu1/aes_top_i/n1210 , \oc8051_xiommu1/aes_top_i/n1211 , 
        \oc8051_xiommu1/aes_top_i/n1212 , \oc8051_xiommu1/aes_top_i/n1213 , 
        \oc8051_xiommu1/aes_top_i/n1214 , \oc8051_xiommu1/aes_top_i/n1215 , 
        \oc8051_xiommu1/aes_top_i/n1216 , \oc8051_xiommu1/aes_top_i/n1217 , 
        \oc8051_xiommu1/aes_top_i/n1218 , \oc8051_xiommu1/aes_top_i/n1219 , 
        \oc8051_xiommu1/aes_top_i/n1220 , \oc8051_xiommu1/aes_top_i/n1221 , 
        \oc8051_xiommu1/aes_top_i/n1222 , \oc8051_xiommu1/aes_top_i/n1223 , 
        \oc8051_xiommu1/aes_top_i/n1224 , \oc8051_xiommu1/aes_top_i/n1225 , 
        \oc8051_xiommu1/aes_top_i/n1226 , \oc8051_xiommu1/aes_top_i/n1227 , 
        \oc8051_xiommu1/aes_top_i/n1228 , \oc8051_xiommu1/aes_top_i/n1229 , 
        \oc8051_xiommu1/aes_top_i/n1230 , \oc8051_xiommu1/aes_top_i/n1231 , 
        \oc8051_xiommu1/aes_top_i/n1232 , \oc8051_xiommu1/aes_top_i/n1233 , 
        \oc8051_xiommu1/aes_top_i/n1234 , \oc8051_xiommu1/aes_top_i/n1235 , 
        \oc8051_xiommu1/aes_top_i/n1236 , \oc8051_xiommu1/aes_top_i/n1237 , 
        \oc8051_xiommu1/aes_top_i/n1238 , \oc8051_xiommu1/aes_top_i/n1239 , 
        \oc8051_xiommu1/aes_top_i/n1240 , \oc8051_xiommu1/aes_top_i/n1241 , 
        \oc8051_xiommu1/aes_top_i/n1242 , \oc8051_xiommu1/aes_top_i/n1243 , 
        \oc8051_xiommu1/aes_top_i/n1244 , \oc8051_xiommu1/aes_top_i/n1245 , 
        \oc8051_xiommu1/aes_top_i/n1246 , \oc8051_xiommu1/aes_top_i/n1247 , 
        \oc8051_xiommu1/aes_top_i/n1248 , \oc8051_xiommu1/aes_top_i/n1249 , 
        \oc8051_xiommu1/aes_top_i/n1250 , \oc8051_xiommu1/aes_top_i/n1251 , 
        \oc8051_xiommu1/aes_top_i/n1252 , \oc8051_xiommu1/aes_top_i/n1253 , 
        \oc8051_xiommu1/aes_top_i/n1254 , \oc8051_xiommu1/aes_top_i/n1255 , 
        \oc8051_xiommu1/aes_top_i/n1256 , \oc8051_xiommu1/aes_top_i/n1257 , 
        \oc8051_xiommu1/aes_top_i/n1258 , \oc8051_xiommu1/aes_top_i/n1259 , 
        \oc8051_xiommu1/aes_top_i/n1260 , \oc8051_xiommu1/aes_top_i/n1261 , 
        \oc8051_xiommu1/aes_top_i/n1262 , \oc8051_xiommu1/aes_top_i/n1263 , 
        \oc8051_xiommu1/aes_top_i/n1264 , \oc8051_xiommu1/aes_top_i/n1265 , 
        \oc8051_xiommu1/aes_top_i/n1266 , \oc8051_xiommu1/aes_top_i/n1267 , 
        \oc8051_xiommu1/aes_top_i/n1268 , \oc8051_xiommu1/aes_top_i/n1269 , 
        \oc8051_xiommu1/aes_top_i/n1270 , \oc8051_xiommu1/aes_top_i/n1271 , 
        \oc8051_xiommu1/aes_top_i/n1272 , \oc8051_xiommu1/aes_top_i/n1273 , 
        \oc8051_xiommu1/aes_top_i/n1274 , \oc8051_xiommu1/aes_top_i/n1275 , 
        \oc8051_xiommu1/aes_top_i/n1276 , \oc8051_xiommu1/aes_top_i/n1277 , 
        \oc8051_xiommu1/aes_top_i/n1278 , \oc8051_xiommu1/aes_top_i/n1279 , 
        \oc8051_xiommu1/aes_top_i/n1280 , \oc8051_xiommu1/aes_top_i/n1281 , 
        \oc8051_xiommu1/aes_top_i/n1282 , \oc8051_xiommu1/aes_top_i/n1283 , 
        \oc8051_xiommu1/aes_top_i/n1284 , \oc8051_xiommu1/aes_top_i/n1285 , 
        \oc8051_xiommu1/aes_top_i/n1286 , \oc8051_xiommu1/aes_top_i/n1287 , 
        \oc8051_xiommu1/aes_top_i/n1288 , \oc8051_xiommu1/aes_top_i/n1289 , 
        \oc8051_xiommu1/aes_top_i/n1290 , \oc8051_xiommu1/aes_top_i/n1291 , 
        \oc8051_xiommu1/aes_top_i/n1292 , \oc8051_xiommu1/aes_top_i/n1293 , 
        \oc8051_xiommu1/aes_top_i/n1294 , \oc8051_xiommu1/aes_top_i/n1295 , 
        \oc8051_xiommu1/aes_top_i/n1296 , \oc8051_xiommu1/aes_top_i/n1297 , 
        \oc8051_xiommu1/aes_top_i/n1298 , \oc8051_xiommu1/aes_top_i/n1299 , 
        \oc8051_xiommu1/aes_top_i/n1300 , \oc8051_xiommu1/aes_top_i/n1301 , 
        \oc8051_xiommu1/aes_top_i/n1302 , \oc8051_xiommu1/aes_top_i/n1303 , 
        \oc8051_xiommu1/aes_top_i/n1304 , \oc8051_xiommu1/aes_top_i/n1305 , 
        \oc8051_xiommu1/aes_top_i/n1306 , \oc8051_xiommu1/aes_top_i/n1307 , 
        \oc8051_xiommu1/aes_top_i/n1308 , \oc8051_xiommu1/aes_top_i/n1309 , 
        \oc8051_xiommu1/aes_top_i/n1310 , \oc8051_xiommu1/aes_top_i/n1311 , 
        \oc8051_xiommu1/aes_top_i/n1312 , \oc8051_xiommu1/aes_top_i/n1313 , 
        \oc8051_xiommu1/aes_top_i/n1314 , \oc8051_xiommu1/aes_top_i/n1315 , 
        \oc8051_xiommu1/aes_top_i/n1316 , \oc8051_xiommu1/aes_top_i/n1317 , 
        \oc8051_xiommu1/aes_top_i/n1318 , \oc8051_xiommu1/aes_top_i/n1319 , 
        \oc8051_xiommu1/aes_top_i/n1320 , \oc8051_xiommu1/aes_top_i/n1321 , 
        \oc8051_xiommu1/aes_top_i/n1322 , \oc8051_xiommu1/aes_top_i/n1323 , 
        \oc8051_xiommu1/aes_top_i/n1324 , \oc8051_xiommu1/aes_top_i/n1325 , 
        \oc8051_xiommu1/aes_top_i/n1326 , \oc8051_xiommu1/aes_top_i/n1327 , 
        \oc8051_xiommu1/aes_top_i/n1328 , \oc8051_xiommu1/aes_top_i/n1329 , 
        \oc8051_xiommu1/aes_top_i/n1330 , \oc8051_xiommu1/aes_top_i/n1331 , 
        \oc8051_xiommu1/aes_top_i/n1332 , \oc8051_xiommu1/aes_top_i/n1333 , 
        \oc8051_xiommu1/aes_top_i/n1334 , \oc8051_xiommu1/aes_top_i/n1335 , 
        \oc8051_xiommu1/aes_top_i/n1336 , \oc8051_xiommu1/aes_top_i/n1337 , 
        \oc8051_xiommu1/aes_top_i/n1338 , \oc8051_xiommu1/aes_top_i/n1339 , 
        \oc8051_xiommu1/aes_top_i/n1340 , \oc8051_xiommu1/aes_top_i/n1341 , 
        \oc8051_xiommu1/aes_top_i/n1342 , \oc8051_xiommu1/aes_top_i/n1343 , 
        \oc8051_xiommu1/aes_top_i/n1344 , \oc8051_xiommu1/aes_top_i/n1345 , 
        \oc8051_xiommu1/aes_top_i/n1346 , \oc8051_xiommu1/aes_top_i/n1347 , 
        \oc8051_xiommu1/aes_top_i/n1348 , \oc8051_xiommu1/aes_top_i/n1349 , 
        \oc8051_xiommu1/aes_top_i/n1350 , \oc8051_xiommu1/aes_top_i/n1351 , 
        \oc8051_xiommu1/aes_top_i/n1352 , \oc8051_xiommu1/aes_top_i/n1353 , 
        \oc8051_xiommu1/aes_top_i/n1354 , \oc8051_xiommu1/aes_top_i/n1355 , 
        \oc8051_xiommu1/aes_top_i/n1356 , \oc8051_xiommu1/aes_top_i/n1357 , 
        \oc8051_xiommu1/aes_top_i/n1358 , \oc8051_xiommu1/aes_top_i/n1359 , 
        \oc8051_xiommu1/aes_top_i/n1360 , \oc8051_xiommu1/aes_top_i/n1361 , 
        \oc8051_xiommu1/aes_top_i/n1362 , \oc8051_xiommu1/aes_top_i/n1363 , 
        \oc8051_xiommu1/aes_top_i/n1364 , \oc8051_xiommu1/aes_top_i/n1365 , 
        \oc8051_xiommu1/aes_top_i/n1366 , \oc8051_xiommu1/aes_top_i/n1367 , 
        \oc8051_xiommu1/aes_top_i/n1368 , \oc8051_xiommu1/aes_top_i/n1369 , 
        \oc8051_xiommu1/aes_top_i/n1370 , \oc8051_xiommu1/aes_top_i/n1371 , 
        \oc8051_xiommu1/aes_top_i/n1372 , \oc8051_xiommu1/aes_top_i/n1373 , 
        \oc8051_xiommu1/aes_top_i/n1374 , \oc8051_xiommu1/aes_top_i/n1375 , 
        \oc8051_xiommu1/aes_top_i/n1376 , \oc8051_xiommu1/aes_top_i/n1377 , 
        \oc8051_xiommu1/aes_top_i/n1378 , \oc8051_xiommu1/aes_top_i/n1379 , 
        \oc8051_xiommu1/aes_top_i/n1380 , \oc8051_xiommu1/aes_top_i/n1381 , 
        \oc8051_xiommu1/aes_top_i/n1382 , \oc8051_xiommu1/aes_top_i/n1383 , 
        \oc8051_xiommu1/aes_top_i/n1384 , \oc8051_xiommu1/aes_top_i/n1385 , 
        \oc8051_xiommu1/aes_top_i/n1386 , \oc8051_xiommu1/aes_top_i/n1387 , 
        \oc8051_xiommu1/aes_top_i/n1388 , \oc8051_xiommu1/aes_top_i/n1389 , 
        \oc8051_xiommu1/aes_top_i/n1390 , \oc8051_xiommu1/aes_top_i/n1391 , 
        \oc8051_xiommu1/aes_top_i/n1392 , \oc8051_xiommu1/aes_top_i/n1393 , 
        \oc8051_xiommu1/aes_top_i/n1394 , \oc8051_xiommu1/aes_top_i/n1395 , 
        \oc8051_xiommu1/aes_top_i/n1396 , \oc8051_xiommu1/aes_top_i/n1397 , 
        \oc8051_xiommu1/aes_top_i/n1398 , \oc8051_xiommu1/aes_top_i/n1399 , 
        \oc8051_xiommu1/aes_top_i/n1400 , \oc8051_xiommu1/aes_top_i/n1401 , 
        \oc8051_xiommu1/aes_top_i/n1402 , \oc8051_xiommu1/aes_top_i/n1403 , 
        \oc8051_xiommu1/aes_top_i/n1404 , \oc8051_xiommu1/aes_top_i/n1405 , 
        \oc8051_xiommu1/aes_top_i/n1406 , \oc8051_xiommu1/aes_top_i/n1407 , 
        \oc8051_xiommu1/aes_top_i/n1408 , \oc8051_xiommu1/aes_top_i/n1409 , 
        \oc8051_xiommu1/aes_top_i/n1410 , \oc8051_xiommu1/aes_top_i/n1411 , 
        \oc8051_xiommu1/aes_top_i/n1412 , \oc8051_xiommu1/aes_top_i/n1413 , 
        \oc8051_xiommu1/aes_top_i/n1414 , \oc8051_xiommu1/aes_top_i/n1415 , 
        \oc8051_xiommu1/aes_top_i/n1416 , \oc8051_xiommu1/aes_top_i/n1417 , 
        \oc8051_xiommu1/aes_top_i/n1418 , \oc8051_xiommu1/aes_top_i/n1419 , 
        \oc8051_xiommu1/aes_top_i/n1420 , \oc8051_xiommu1/aes_top_i/n1421 , 
        \oc8051_xiommu1/aes_top_i/n1422 , \oc8051_xiommu1/aes_top_i/n1423 , 
        \oc8051_xiommu1/aes_top_i/n1424 , \oc8051_xiommu1/aes_top_i/n1425 , 
        \oc8051_xiommu1/aes_top_i/n1426 , \oc8051_xiommu1/aes_top_i/n1427 , 
        \oc8051_xiommu1/aes_top_i/n1428 , \oc8051_xiommu1/aes_top_i/n1429 , 
        \oc8051_xiommu1/aes_top_i/n1430 , \oc8051_xiommu1/aes_top_i/n1431 , 
        \oc8051_xiommu1/aes_top_i/n1432 , \oc8051_xiommu1/aes_top_i/n1433 , 
        \oc8051_xiommu1/aes_top_i/n1434 , \oc8051_xiommu1/aes_top_i/n1435 , 
        \oc8051_xiommu1/aes_top_i/n1436 , \oc8051_xiommu1/aes_top_i/n1437 , 
        \oc8051_xiommu1/aes_top_i/n1438 , \oc8051_xiommu1/aes_top_i/n1439 , 
        \oc8051_xiommu1/aes_top_i/n1440 , \oc8051_xiommu1/aes_top_i/n1441 , 
        \oc8051_xiommu1/aes_top_i/n1442 , \oc8051_xiommu1/aes_top_i/n1443 , 
        \oc8051_xiommu1/aes_top_i/n1444 , \oc8051_xiommu1/aes_top_i/n1445 , 
        \oc8051_xiommu1/aes_top_i/n1446 , \oc8051_xiommu1/aes_top_i/n1447 , 
        \oc8051_xiommu1/aes_top_i/n1448 , \oc8051_xiommu1/aes_top_i/n1449 , 
        \oc8051_xiommu1/aes_top_i/n1450 , \oc8051_xiommu1/aes_top_i/n1451 , 
        \oc8051_xiommu1/aes_top_i/n1452 , \oc8051_xiommu1/aes_top_i/n1453 , 
        \oc8051_xiommu1/aes_top_i/n1454 , \oc8051_xiommu1/aes_top_i/n1455 , 
        \oc8051_xiommu1/aes_top_i/n1456 , \oc8051_xiommu1/aes_top_i/n1457 , 
        \oc8051_xiommu1/aes_top_i/n1458 , \oc8051_xiommu1/aes_top_i/n1459 , 
        \oc8051_xiommu1/aes_top_i/n1460 , \oc8051_xiommu1/aes_top_i/n1461 , 
        \oc8051_xiommu1/aes_top_i/n1462 , \oc8051_xiommu1/aes_top_i/n1463 , 
        \oc8051_xiommu1/aes_top_i/n1464 , \oc8051_xiommu1/aes_top_i/n1465 , 
        \oc8051_xiommu1/aes_top_i/n1466 , \oc8051_xiommu1/aes_top_i/n1467 , 
        \oc8051_xiommu1/aes_top_i/n1468 , \oc8051_xiommu1/aes_top_i/n1469 , 
        \oc8051_xiommu1/aes_top_i/n1470 , \oc8051_xiommu1/aes_top_i/n1471 , 
        \oc8051_xiommu1/aes_top_i/n1472 , \oc8051_xiommu1/aes_top_i/n1473 , 
        \oc8051_xiommu1/aes_top_i/n1474 , \oc8051_xiommu1/aes_top_i/n1475 , 
        \oc8051_xiommu1/aes_top_i/n1476 , \oc8051_xiommu1/aes_top_i/n1477 , 
        \oc8051_xiommu1/aes_top_i/n1478 , \oc8051_xiommu1/aes_top_i/n1479 , 
        \oc8051_xiommu1/aes_top_i/n1480 , \oc8051_xiommu1/aes_top_i/n1481 , 
        \oc8051_xiommu1/aes_top_i/n1482 , \oc8051_xiommu1/aes_top_i/n1483 , 
        \oc8051_xiommu1/aes_top_i/n1484 , \oc8051_xiommu1/aes_top_i/n1485 , 
        \oc8051_xiommu1/aes_top_i/n1486 , \oc8051_xiommu1/aes_top_i/n1487 , 
        \oc8051_xiommu1/aes_top_i/n1488 , \oc8051_xiommu1/aes_top_i/n1489 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n70 , \oc8051_xiommu1/oc8051_procarbiter_i/n71 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n72 , \oc8051_xiommu1/oc8051_procarbiter_i/n78 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n79 , \oc8051_xiommu1/oc8051_memarbiter_i/n48 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n49 , \oc8051_xiommu1/oc8051_memarbiter_i/n50 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n51 , \oc8051_xiommu1/oc8051_memarbiter_i/n52 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n53 , \oc8051_xiommu1/oc8051_memarbiter_i/n54 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n55 , \oc8051_xiommu1/oc8051_memarbiter_i/n56 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n57 , \oc8051_xiommu1/oc8051_memarbiter_i/n58 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n59 , \oc8051_xiommu1/oc8051_memarbiter_i/n60 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n61 , \oc8051_xiommu1/oc8051_memarbiter_i/n62 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n63 , \oc8051_xiommu1/oc8051_memarbiter_i/n64 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n65 , \oc8051_xiommu1/oc8051_memarbiter_i/n66 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n67 , \oc8051_xiommu1/oc8051_memarbiter_i/n68 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n69 , \oc8051_xiommu1/oc8051_memarbiter_i/n70 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n71 , \oc8051_xiommu1/oc8051_memarbiter_i/n72 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n73 , \oc8051_xiommu1/oc8051_memarbiter_i/n74 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n75 , \oc8051_xiommu1/oc8051_memarbiter_i/n76 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n77 , \oc8051_xiommu1/oc8051_memarbiter_i/n78 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n79 , \oc8051_xiommu1/oc8051_memarbiter_i/n80 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n81 , \oc8051_xiommu1/oc8051_memarbiter_i/n82 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n83 , \oc8051_xiommu1/oc8051_memarbiter_i/n108 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n109 , \oc8051_xiommu1/oc8051_memarbiter_i/n110 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n111 , \oc8051_xiommu1/oc8051_memarbiter_i/n112 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n113 , \oc8051_xiommu1/oc8051_memarbiter_i/n114 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n115 , \oc8051_xiommu1/oc8051_memarbiter_i/n116 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n117 , \oc8051_xiommu1/oc8051_memarbiter_i/n118 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n119 , \oc8051_xiommu1/oc8051_memarbiter_i/n120 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n121 , \oc8051_xiommu1/oc8051_memarbiter_i/n122 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n123 , \oc8051_xiommu1/oc8051_memarbiter_i/n124 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n125 , \oc8051_xiommu1/oc8051_memarbiter_i/n126 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n127 , \oc8051_xiommu1/oc8051_memarbiter_i/n128 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n129 , \oc8051_xiommu1/oc8051_memarbiter_i/n130 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n131 , \oc8051_xiommu1/oc8051_memarbiter_i/n152 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n156 , \oc8051_xiommu1/oc8051_memarbiter_i/n157 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n158 , \oc8051_xiommu1/oc8051_memarbiter_i/n159 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n168 , \oc8051_xiommu1/oc8051_memarbiter_i/n169 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n170 , \oc8051_xiommu1/oc8051_memarbiter_i/n171 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n172 , \oc8051_xiommu1/oc8051_memarbiter_i/n173 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n174 , \oc8051_xiommu1/oc8051_memarbiter_i/n187 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n188 , \oc8051_xiommu1/oc8051_memarbiter_i/n189 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n190 , \oc8051_xiommu1/oc8051_memarbiter_i/n201 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n202 , \oc8051_xiommu1/oc8051_memarbiter_i/n203 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n204 , \oc8051_xiommu1/oc8051_page_table_i/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/n5 , \oc8051_xiommu1/oc8051_page_table_i/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/n8 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 , \oc8051_xiommu1/oc8051_page_table_i/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/n34 , \oc8051_xiommu1/oc8051_page_table_i/n59 , 
        \oc8051_xiommu1/oc8051_page_table_i/n84 , \oc8051_xiommu1/oc8051_page_table_i/n85 , 
        \oc8051_xiommu1/oc8051_page_table_i/n86 , \oc8051_xiommu1/oc8051_page_table_i/n87 , 
        \oc8051_xiommu1/oc8051_page_table_i/n89 , \oc8051_xiommu1/oc8051_page_table_i/n93 , 
        \oc8051_xiommu1/oc8051_page_table_i/n94 , \oc8051_xiommu1/oc8051_page_table_i/n95 , 
        \oc8051_xiommu1/oc8051_page_table_i/n96 , \oc8051_xiommu1/oc8051_page_table_i/n97 , 
        \oc8051_xiommu1/oc8051_page_table_i/n98 , \oc8051_xiommu1/oc8051_page_table_i/n99 , 
        \oc8051_xiommu1/oc8051_page_table_i/n100 , \oc8051_xiommu1/oc8051_page_table_i/n109 , 
        \oc8051_xiommu1/oc8051_page_table_i/n110 , \oc8051_xiommu1/oc8051_page_table_i/n111 , 
        \oc8051_xiommu1/oc8051_page_table_i/n112 , \oc8051_xiommu1/oc8051_page_table_i/n113 , 
        \oc8051_xiommu1/oc8051_page_table_i/n114 , \oc8051_xiommu1/oc8051_page_table_i/n115 , 
        \oc8051_xiommu1/oc8051_page_table_i/n116 , \oc8051_xiommu1/oc8051_page_table_i/n118 , 
        \oc8051_xiommu1/oc8051_page_table_i/n119 , \oc8051_xiommu1/oc8051_page_table_i/n120 , 
        \oc8051_xiommu1/oc8051_page_table_i/n121 , \oc8051_xiommu1/oc8051_page_table_i/n122 , 
        \oc8051_xiommu1/oc8051_page_table_i/n123 , \oc8051_xiommu1/oc8051_page_table_i/n124 , 
        \oc8051_xiommu1/oc8051_page_table_i/n125 , \oc8051_xiommu1/oc8051_page_table_i/n128 , 
        \oc8051_xiommu1/oc8051_page_table_i/n129 , \oc8051_xiommu1/oc8051_page_table_i/n130 , 
        \oc8051_xiommu1/oc8051_page_table_i/n131 , \oc8051_xiommu1/oc8051_page_table_i/n132 , 
        \oc8051_xiommu1/oc8051_page_table_i/n133 , \oc8051_xiommu1/oc8051_page_table_i/n134 , 
        \oc8051_xiommu1/oc8051_page_table_i/n135 , \oc8051_xiommu1/oc8051_page_table_i/n144 , 
        \oc8051_xiommu1/oc8051_page_table_i/n145 , \oc8051_xiommu1/oc8051_page_table_i/n146 , 
        \oc8051_xiommu1/oc8051_page_table_i/n147 , \oc8051_xiommu1/oc8051_page_table_i/n148 , 
        \oc8051_xiommu1/oc8051_page_table_i/n149 , \oc8051_xiommu1/oc8051_page_table_i/n150 , 
        \oc8051_xiommu1/oc8051_page_table_i/n151 , \oc8051_xiommu1/oc8051_page_table_i/n194 , 
        \oc8051_xiommu1/oc8051_page_table_i/n195 , \oc8051_xiommu1/oc8051_page_table_i/n196 , 
        \oc8051_xiommu1/oc8051_page_table_i/n197 , \oc8051_xiommu1/oc8051_page_table_i/n198 , 
        \oc8051_xiommu1/oc8051_page_table_i/n199 , \oc8051_xiommu1/oc8051_page_table_i/n200 , 
        \oc8051_xiommu1/oc8051_page_table_i/n201 , \oc8051_xiommu1/oc8051_page_table_i/n202 , 
        \oc8051_xiommu1/oc8051_page_table_i/n203 , \oc8051_xiommu1/oc8051_page_table_i/n204 , 
        \oc8051_xiommu1/oc8051_page_table_i/n205 , \oc8051_xiommu1/oc8051_page_table_i/n206 , 
        \oc8051_xiommu1/oc8051_page_table_i/n207 , \oc8051_xiommu1/oc8051_page_table_i/n208 , 
        \oc8051_xiommu1/oc8051_page_table_i/n209 , \oc8051_xiommu1/oc8051_page_table_i/n210 , 
        \oc8051_xiommu1/oc8051_page_table_i/n211 , \oc8051_xiommu1/oc8051_page_table_i/n212 , 
        \oc8051_xiommu1/oc8051_page_table_i/n213 , \oc8051_xiommu1/oc8051_page_table_i/n214 , 
        \oc8051_xiommu1/oc8051_page_table_i/n215 , \oc8051_xiommu1/oc8051_page_table_i/n216 , 
        \oc8051_xiommu1/oc8051_page_table_i/n217 , \oc8051_xiommu1/oc8051_page_table_i/n218 , 
        \oc8051_xiommu1/oc8051_page_table_i/n219 , \oc8051_xiommu1/oc8051_page_table_i/n220 , 
        \oc8051_xiommu1/oc8051_page_table_i/n221 , \oc8051_xiommu1/oc8051_page_table_i/n222 , 
        \oc8051_xiommu1/oc8051_page_table_i/n223 , \oc8051_xiommu1/oc8051_page_table_i/n224 , 
        \oc8051_xiommu1/oc8051_page_table_i/n225 , \oc8051_xiommu1/oc8051_page_table_i/n226 , 
        \oc8051_xiommu1/oc8051_page_table_i/n227 , \oc8051_xiommu1/oc8051_page_table_i/n228 , 
        \oc8051_xiommu1/oc8051_page_table_i/n229 , \oc8051_xiommu1/oc8051_page_table_i/n230 , 
        \oc8051_xiommu1/oc8051_page_table_i/n231 , \oc8051_xiommu1/oc8051_page_table_i/n232 , 
        \oc8051_xiommu1/oc8051_page_table_i/n233 , \oc8051_xiommu1/oc8051_page_table_i/n234 , 
        \oc8051_xiommu1/oc8051_page_table_i/n235 , \oc8051_xiommu1/oc8051_page_table_i/n236 , 
        \oc8051_xiommu1/oc8051_page_table_i/n237 , \oc8051_xiommu1/oc8051_page_table_i/n238 , 
        \oc8051_xiommu1/oc8051_page_table_i/n239 , \oc8051_xiommu1/oc8051_page_table_i/n240 , 
        \oc8051_xiommu1/oc8051_page_table_i/n241 , \oc8051_xiommu1/oc8051_page_table_i/n242 , 
        \oc8051_xiommu1/oc8051_page_table_i/n243 , \oc8051_xiommu1/oc8051_page_table_i/n244 , 
        \oc8051_xiommu1/oc8051_page_table_i/n245 , \oc8051_xiommu1/oc8051_page_table_i/n246 , 
        \oc8051_xiommu1/oc8051_page_table_i/n247 , \oc8051_xiommu1/oc8051_page_table_i/n248 , 
        \oc8051_xiommu1/oc8051_page_table_i/n249 , \oc8051_xiommu1/oc8051_page_table_i/n250 , 
        \oc8051_xiommu1/oc8051_page_table_i/n251 , \oc8051_xiommu1/oc8051_page_table_i/n252 , 
        \oc8051_xiommu1/oc8051_page_table_i/n253 , \oc8051_xiommu1/oc8051_page_table_i/n254 , 
        \oc8051_xiommu1/oc8051_page_table_i/n255 , \oc8051_xiommu1/oc8051_page_table_i/n256 , 
        \oc8051_xiommu1/oc8051_page_table_i/n257 , \oc8051_xiommu1/oc8051_page_table_i/n258 , 
        \oc8051_xiommu1/oc8051_page_table_i/n259 , \oc8051_xiommu1/oc8051_page_table_i/n260 , 
        \oc8051_xiommu1/oc8051_page_table_i/n261 , \oc8051_xiommu1/oc8051_page_table_i/n262 , 
        \oc8051_xiommu1/oc8051_page_table_i/n263 , \oc8051_xiommu1/oc8051_page_table_i/n264 , 
        \oc8051_xiommu1/oc8051_page_table_i/n265 , \oc8051_xiommu1/oc8051_page_table_i/n266 , 
        \oc8051_xiommu1/oc8051_page_table_i/n267 , \oc8051_xiommu1/oc8051_page_table_i/n268 , 
        \oc8051_xiommu1/oc8051_page_table_i/n269 , \oc8051_xiommu1/oc8051_page_table_i/n270 , 
        \oc8051_xiommu1/oc8051_page_table_i/n271 , \oc8051_xiommu1/oc8051_page_table_i/n272 , 
        \oc8051_xiommu1/oc8051_page_table_i/n273 , \oc8051_xiommu1/oc8051_page_table_i/n274 , 
        \oc8051_xiommu1/oc8051_page_table_i/n275 , \oc8051_xiommu1/oc8051_page_table_i/n276 , 
        \oc8051_xiommu1/oc8051_page_table_i/n277 , \oc8051_xiommu1/oc8051_page_table_i/n278 , 
        \oc8051_xiommu1/oc8051_page_table_i/n279 , \oc8051_xiommu1/oc8051_page_table_i/n280 , 
        \oc8051_xiommu1/oc8051_page_table_i/n281 , \oc8051_xiommu1/oc8051_page_table_i/n282 , 
        \oc8051_xiommu1/oc8051_page_table_i/n283 , \oc8051_xiommu1/oc8051_page_table_i/n284 , 
        \oc8051_xiommu1/oc8051_page_table_i/n285 , \oc8051_xiommu1/oc8051_page_table_i/n286 , 
        \oc8051_xiommu1/oc8051_page_table_i/n287 , \oc8051_xiommu1/oc8051_page_table_i/n288 , 
        \oc8051_xiommu1/oc8051_page_table_i/n289 , \oc8051_xiommu1/oc8051_page_table_i/n290 , 
        \oc8051_xiommu1/oc8051_page_table_i/n291 , \oc8051_xiommu1/oc8051_page_table_i/n292 , 
        \oc8051_xiommu1/oc8051_page_table_i/n293 , \oc8051_xiommu1/oc8051_page_table_i/n294 , 
        \oc8051_xiommu1/oc8051_page_table_i/n295 , \oc8051_xiommu1/oc8051_page_table_i/n296 , 
        \oc8051_xiommu1/oc8051_page_table_i/n297 , \oc8051_xiommu1/oc8051_page_table_i/n298 , 
        \oc8051_xiommu1/oc8051_page_table_i/n299 , \oc8051_xiommu1/oc8051_page_table_i/n300 , 
        \oc8051_xiommu1/oc8051_page_table_i/n301 , \oc8051_xiommu1/oc8051_page_table_i/n302 , 
        \oc8051_xiommu1/oc8051_page_table_i/n303 , \oc8051_xiommu1/oc8051_page_table_i/n304 , 
        \oc8051_xiommu1/oc8051_page_table_i/n305 , \oc8051_xiommu1/oc8051_page_table_i/n306 , 
        \oc8051_xiommu1/oc8051_page_table_i/n307 , \oc8051_xiommu1/oc8051_page_table_i/n308 , 
        \oc8051_xiommu1/oc8051_page_table_i/n309 , \oc8051_xiommu1/oc8051_page_table_i/n310 , 
        \oc8051_xiommu1/oc8051_page_table_i/n311 , \oc8051_xiommu1/oc8051_page_table_i/n312 , 
        \oc8051_xiommu1/oc8051_page_table_i/n313 , \oc8051_xiommu1/oc8051_page_table_i/n314 , 
        \oc8051_xiommu1/oc8051_page_table_i/n315 , \oc8051_xiommu1/oc8051_page_table_i/n316 , 
        \oc8051_xiommu1/oc8051_page_table_i/n317 , \oc8051_xiommu1/oc8051_page_table_i/n318 , 
        \oc8051_xiommu1/oc8051_page_table_i/n319 , \oc8051_xiommu1/oc8051_page_table_i/n320 , 
        \oc8051_xiommu1/oc8051_page_table_i/n321 , \oc8051_xiommu1/oc8051_page_table_i/n322 , 
        \oc8051_xiommu1/oc8051_page_table_i/n323 , \oc8051_xiommu1/oc8051_page_table_i/n324 , 
        \oc8051_xiommu1/oc8051_page_table_i/n325 , \oc8051_xiommu1/oc8051_page_table_i/n326 , 
        \oc8051_xiommu1/oc8051_page_table_i/n327 , \oc8051_xiommu1/oc8051_page_table_i/n328 , 
        \oc8051_xiommu1/oc8051_page_table_i/n329 , \oc8051_xiommu1/oc8051_page_table_i/n330 , 
        \oc8051_xiommu1/oc8051_page_table_i/n331 , \oc8051_xiommu1/oc8051_page_table_i/n332 , 
        \oc8051_xiommu1/oc8051_page_table_i/n333 , \oc8051_xiommu1/oc8051_page_table_i/n334 , 
        \oc8051_xiommu1/oc8051_page_table_i/n335 , \oc8051_xiommu1/oc8051_page_table_i/n336 , 
        \oc8051_xiommu1/oc8051_page_table_i/n337 , \oc8051_xiommu1/oc8051_page_table_i/n338 , 
        \oc8051_xiommu1/oc8051_page_table_i/n339 , \oc8051_xiommu1/oc8051_page_table_i/n340 , 
        \oc8051_xiommu1/oc8051_page_table_i/n341 , \oc8051_xiommu1/oc8051_page_table_i/n342 , 
        \oc8051_xiommu1/oc8051_page_table_i/n343 , \oc8051_xiommu1/oc8051_page_table_i/n344 , 
        \oc8051_xiommu1/oc8051_page_table_i/n345 , \oc8051_xiommu1/oc8051_page_table_i/n346 , 
        \oc8051_xiommu1/oc8051_page_table_i/n347 , \oc8051_xiommu1/oc8051_page_table_i/n348 , 
        \oc8051_xiommu1/oc8051_page_table_i/n349 , \oc8051_xiommu1/oc8051_page_table_i/n350 , 
        \oc8051_xiommu1/oc8051_page_table_i/n351 , \oc8051_xiommu1/oc8051_page_table_i/n352 , 
        \oc8051_xiommu1/oc8051_page_table_i/n353 , \oc8051_xiommu1/oc8051_page_table_i/n354 , 
        \oc8051_xiommu1/oc8051_page_table_i/n355 , \oc8051_xiommu1/oc8051_page_table_i/n356 , 
        \oc8051_xiommu1/oc8051_page_table_i/n357 , \oc8051_xiommu1/oc8051_page_table_i/n358 , 
        \oc8051_xiommu1/oc8051_page_table_i/n359 , \oc8051_xiommu1/oc8051_page_table_i/n360 , 
        \oc8051_xiommu1/oc8051_page_table_i/n361 , \oc8051_xiommu1/oc8051_page_table_i/n362 , 
        \oc8051_xiommu1/oc8051_page_table_i/n363 , \oc8051_xiommu1/oc8051_page_table_i/n364 , 
        \oc8051_xiommu1/oc8051_page_table_i/n365 , \oc8051_xiommu1/oc8051_page_table_i/n366 , 
        \oc8051_xiommu1/oc8051_page_table_i/n367 , \oc8051_xiommu1/oc8051_page_table_i/n368 , 
        \oc8051_xiommu1/oc8051_page_table_i/n369 , \oc8051_xiommu1/oc8051_page_table_i/n370 , 
        \oc8051_xiommu1/oc8051_page_table_i/n371 , \oc8051_xiommu1/oc8051_page_table_i/n372 , 
        \oc8051_xiommu1/oc8051_page_table_i/n373 , \oc8051_xiommu1/oc8051_page_table_i/n374 , 
        \oc8051_xiommu1/oc8051_page_table_i/n375 , \oc8051_xiommu1/oc8051_page_table_i/n376 , 
        \oc8051_xiommu1/oc8051_page_table_i/n377 , \oc8051_xiommu1/oc8051_page_table_i/n378 , 
        \oc8051_xiommu1/oc8051_page_table_i/n379 , \oc8051_xiommu1/oc8051_page_table_i/n380 , 
        \oc8051_xiommu1/oc8051_page_table_i/n381 , \oc8051_xiommu1/oc8051_page_table_i/n382 , 
        \oc8051_xiommu1/oc8051_page_table_i/n383 , \oc8051_xiommu1/oc8051_page_table_i/n384 , 
        \oc8051_xiommu1/oc8051_page_table_i/n385 , \oc8051_xiommu1/oc8051_page_table_i/n386 , 
        \oc8051_xiommu1/oc8051_page_table_i/n387 , \oc8051_xiommu1/oc8051_page_table_i/n388 , 
        \oc8051_xiommu1/oc8051_page_table_i/n389 , \oc8051_xiommu1/oc8051_page_table_i/n390 , 
        \oc8051_xiommu1/oc8051_page_table_i/n391 , \oc8051_xiommu1/oc8051_page_table_i/n392 , 
        \oc8051_xiommu1/oc8051_page_table_i/n393 , \oc8051_xiommu1/oc8051_page_table_i/n394 , 
        \oc8051_xiommu1/oc8051_page_table_i/n395 , \oc8051_xiommu1/oc8051_page_table_i/n396 , 
        \oc8051_xiommu1/oc8051_page_table_i/n397 , \oc8051_xiommu1/oc8051_page_table_i/n398 , 
        \oc8051_xiommu1/oc8051_page_table_i/n399 , \oc8051_xiommu1/oc8051_page_table_i/n400 , 
        \oc8051_xiommu1/oc8051_page_table_i/n401 , \oc8051_xiommu1/oc8051_page_table_i/n402 , 
        \oc8051_xiommu1/oc8051_page_table_i/n403 , \oc8051_xiommu1/oc8051_page_table_i/n404 , 
        \oc8051_xiommu1/oc8051_page_table_i/n405 , \oc8051_xiommu1/oc8051_page_table_i/n406 , 
        \oc8051_xiommu1/oc8051_page_table_i/n407 , \oc8051_xiommu1/oc8051_page_table_i/n408 , 
        \oc8051_xiommu1/oc8051_page_table_i/n409 , \oc8051_xiommu1/oc8051_page_table_i/n410 , 
        \oc8051_xiommu1/oc8051_page_table_i/n411 , \oc8051_xiommu1/oc8051_page_table_i/n412 , 
        \oc8051_xiommu1/oc8051_page_table_i/n413 , \oc8051_xiommu1/oc8051_page_table_i/n414 , 
        \oc8051_xiommu1/oc8051_page_table_i/n415 , \oc8051_xiommu1/oc8051_page_table_i/n416 , 
        \oc8051_xiommu1/oc8051_page_table_i/n417 , \oc8051_xiommu1/oc8051_page_table_i/n418 , 
        \oc8051_xiommu1/oc8051_page_table_i/n419 , \oc8051_xiommu1/oc8051_page_table_i/n420 , 
        \oc8051_xiommu1/oc8051_page_table_i/n421 , \oc8051_xiommu1/oc8051_page_table_i/n422 , 
        \oc8051_xiommu1/oc8051_page_table_i/n423 , \oc8051_xiommu1/oc8051_page_table_i/n424 , 
        \oc8051_xiommu1/oc8051_page_table_i/n425 , \oc8051_xiommu1/oc8051_page_table_i/n426 , 
        \oc8051_xiommu1/oc8051_page_table_i/n427 , \oc8051_xiommu1/oc8051_page_table_i/n428 , 
        \oc8051_xiommu1/oc8051_page_table_i/n429 , \oc8051_xiommu1/oc8051_page_table_i/n430 , 
        \oc8051_xiommu1/oc8051_page_table_i/n431 , \oc8051_xiommu1/oc8051_page_table_i/n432 , 
        \oc8051_xiommu1/oc8051_page_table_i/n433 , \oc8051_xiommu1/oc8051_page_table_i/n434 , 
        \oc8051_xiommu1/oc8051_page_table_i/n435 , \oc8051_xiommu1/oc8051_page_table_i/n436 , 
        \oc8051_xiommu1/oc8051_page_table_i/n437 , \oc8051_xiommu1/oc8051_page_table_i/n438 , 
        \oc8051_xiommu1/oc8051_page_table_i/n439 , \oc8051_xiommu1/oc8051_page_table_i/n440 , 
        \oc8051_xiommu1/oc8051_page_table_i/n441 , \oc8051_xiommu1/oc8051_page_table_i/n442 , 
        \oc8051_xiommu1/oc8051_page_table_i/n443 , \oc8051_xiommu1/oc8051_page_table_i/n444 , 
        \oc8051_xiommu1/oc8051_page_table_i/n445 , \oc8051_xiommu1/oc8051_page_table_i/n446 , 
        \oc8051_xiommu1/oc8051_page_table_i/n447 , \oc8051_xiommu1/oc8051_page_table_i/n448 , 
        \oc8051_xiommu1/oc8051_page_table_i/n449 , \oc8051_xiommu1/oc8051_page_table_i/n483 , 
        \oc8051_xiommu1/oc8051_page_table_i/n484 , \oc8051_xiommu1/oc8051_page_table_i/n485 , 
        \oc8051_xiommu1/oc8051_page_table_i/n486 , \oc8051_xiommu1/oc8051_page_table_i/n487 , 
        \oc8051_xiommu1/oc8051_page_table_i/n488 , \oc8051_xiommu1/oc8051_page_table_i/n489 , 
        \oc8051_xiommu1/oc8051_page_table_i/n490 , \oc8051_xiommu1/oc8051_page_table_i/n491 , 
        \oc8051_xiommu1/oc8051_page_table_i/n492 , \oc8051_xiommu1/oc8051_page_table_i/n493 , 
        \oc8051_xiommu1/oc8051_page_table_i/n494 , \oc8051_xiommu1/oc8051_page_table_i/n495 , 
        \oc8051_xiommu1/oc8051_page_table_i/n496 , \oc8051_xiommu1/oc8051_page_table_i/n497 , 
        \oc8051_xiommu1/oc8051_page_table_i/n498 , \oc8051_xiommu1/oc8051_page_table_i/n499 , 
        \oc8051_xiommu1/oc8051_page_table_i/n500 , \oc8051_xiommu1/oc8051_page_table_i/n501 , 
        \oc8051_xiommu1/oc8051_page_table_i/n502 , \oc8051_xiommu1/oc8051_page_table_i/n503 , 
        \oc8051_xiommu1/oc8051_page_table_i/n504 , \oc8051_xiommu1/oc8051_page_table_i/n505 , 
        \oc8051_xiommu1/oc8051_page_table_i/n506 , \oc8051_xiommu1/oc8051_page_table_i/n507 , 
        \oc8051_xiommu1/oc8051_page_table_i/n508 , \oc8051_xiommu1/oc8051_page_table_i/n509 , 
        \oc8051_xiommu1/oc8051_page_table_i/n510 , \oc8051_xiommu1/oc8051_page_table_i/n511 , 
        \oc8051_xiommu1/oc8051_page_table_i/n512 , \oc8051_xiommu1/oc8051_page_table_i/n513 , 
        \oc8051_xiommu1/oc8051_page_table_i/n514 , \oc8051_xiommu1/oc8051_page_table_i/n515 , 
        \oc8051_xiommu1/oc8051_page_table_i/n516 , \oc8051_xiommu1/oc8051_page_table_i/n517 , 
        \oc8051_xiommu1/oc8051_page_table_i/n518 , \oc8051_xiommu1/oc8051_page_table_i/n519 , 
        \oc8051_xiommu1/oc8051_page_table_i/n520 , \oc8051_xiommu1/oc8051_page_table_i/n521 , 
        \oc8051_xiommu1/oc8051_page_table_i/n522 , \oc8051_xiommu1/oc8051_page_table_i/n523 , 
        \oc8051_xiommu1/oc8051_page_table_i/n524 , \oc8051_xiommu1/oc8051_page_table_i/n525 , 
        \oc8051_xiommu1/oc8051_page_table_i/n526 , \oc8051_xiommu1/oc8051_page_table_i/n527 , 
        \oc8051_xiommu1/oc8051_page_table_i/n528 , \oc8051_xiommu1/oc8051_page_table_i/n529 , 
        \oc8051_xiommu1/oc8051_page_table_i/n530 , \oc8051_xiommu1/oc8051_page_table_i/n531 , 
        \oc8051_xiommu1/oc8051_page_table_i/n532 , \oc8051_xiommu1/oc8051_page_table_i/n533 , 
        \oc8051_xiommu1/oc8051_page_table_i/n534 , \oc8051_xiommu1/oc8051_page_table_i/n535 , 
        \oc8051_xiommu1/oc8051_page_table_i/n536 , \oc8051_xiommu1/oc8051_page_table_i/n537 , 
        \oc8051_xiommu1/oc8051_page_table_i/n538 , \oc8051_xiommu1/oc8051_page_table_i/n539 , 
        \oc8051_xiommu1/oc8051_page_table_i/n540 , \oc8051_xiommu1/oc8051_page_table_i/n541 , 
        \oc8051_xiommu1/oc8051_page_table_i/n542 , \oc8051_xiommu1/oc8051_page_table_i/n543 , 
        \oc8051_xiommu1/oc8051_page_table_i/n544 , \oc8051_xiommu1/oc8051_page_table_i/n545 , 
        \oc8051_xiommu1/oc8051_page_table_i/n546 , \oc8051_xiommu1/oc8051_page_table_i/n547 , 
        \oc8051_xiommu1/oc8051_page_table_i/n548 , \oc8051_xiommu1/oc8051_page_table_i/n549 , 
        \oc8051_xiommu1/oc8051_page_table_i/n550 , \oc8051_xiommu1/oc8051_page_table_i/n551 , 
        \oc8051_xiommu1/oc8051_page_table_i/n552 , \oc8051_xiommu1/oc8051_page_table_i/n553 , 
        \oc8051_xiommu1/oc8051_page_table_i/n554 , \oc8051_xiommu1/oc8051_page_table_i/n555 , 
        \oc8051_xiommu1/oc8051_page_table_i/n556 , \oc8051_xiommu1/oc8051_page_table_i/n557 , 
        \oc8051_xiommu1/oc8051_page_table_i/n558 , \oc8051_xiommu1/oc8051_page_table_i/n559 , 
        \oc8051_xiommu1/oc8051_page_table_i/n560 , \oc8051_xiommu1/oc8051_page_table_i/n561 , 
        \oc8051_xiommu1/oc8051_page_table_i/n562 , \oc8051_xiommu1/oc8051_page_table_i/n563 , 
        \oc8051_xiommu1/oc8051_page_table_i/n564 , \oc8051_xiommu1/oc8051_page_table_i/n565 , 
        \oc8051_xiommu1/oc8051_page_table_i/n566 , \oc8051_xiommu1/oc8051_page_table_i/n567 , 
        \oc8051_xiommu1/oc8051_page_table_i/n568 , \oc8051_xiommu1/oc8051_page_table_i/n569 , 
        \oc8051_xiommu1/oc8051_page_table_i/n570 , \oc8051_xiommu1/oc8051_page_table_i/n571 , 
        \oc8051_xiommu1/oc8051_page_table_i/n572 , \oc8051_xiommu1/oc8051_page_table_i/n573 , 
        \oc8051_xiommu1/oc8051_page_table_i/n574 , \oc8051_xiommu1/oc8051_page_table_i/n575 , 
        \oc8051_xiommu1/oc8051_page_table_i/n576 , \oc8051_xiommu1/oc8051_page_table_i/n577 , 
        \oc8051_xiommu1/oc8051_page_table_i/n578 , \oc8051_xiommu1/oc8051_page_table_i/n579 , 
        \oc8051_xiommu1/oc8051_page_table_i/n580 , \oc8051_xiommu1/oc8051_page_table_i/n581 , 
        \oc8051_xiommu1/oc8051_page_table_i/n582 , \oc8051_xiommu1/oc8051_page_table_i/n583 , 
        \oc8051_xiommu1/oc8051_page_table_i/n584 , \oc8051_xiommu1/oc8051_page_table_i/n585 , 
        \oc8051_xiommu1/oc8051_page_table_i/n586 , \oc8051_xiommu1/oc8051_page_table_i/n587 , 
        \oc8051_xiommu1/oc8051_page_table_i/n588 , \oc8051_xiommu1/oc8051_page_table_i/n589 , 
        \oc8051_xiommu1/oc8051_page_table_i/n590 , \oc8051_xiommu1/oc8051_page_table_i/n591 , 
        \oc8051_xiommu1/oc8051_page_table_i/n592 , \oc8051_xiommu1/oc8051_page_table_i/n593 , 
        \oc8051_xiommu1/oc8051_page_table_i/n594 , \oc8051_xiommu1/oc8051_page_table_i/n595 , 
        \oc8051_xiommu1/oc8051_page_table_i/n596 , \oc8051_xiommu1/oc8051_page_table_i/n597 , 
        \oc8051_xiommu1/oc8051_page_table_i/n598 , \oc8051_xiommu1/oc8051_page_table_i/n599 , 
        \oc8051_xiommu1/oc8051_page_table_i/n600 , \oc8051_xiommu1/oc8051_page_table_i/n601 , 
        \oc8051_xiommu1/oc8051_page_table_i/n602 , \oc8051_xiommu1/oc8051_page_table_i/n603 , 
        \oc8051_xiommu1/oc8051_page_table_i/n604 , \oc8051_xiommu1/oc8051_page_table_i/n605 , 
        \oc8051_xiommu1/oc8051_page_table_i/n606 , \oc8051_xiommu1/oc8051_page_table_i/n607 , 
        \oc8051_xiommu1/oc8051_page_table_i/n608 , \oc8051_xiommu1/oc8051_page_table_i/n609 , 
        \oc8051_xiommu1/oc8051_page_table_i/n610 , \oc8051_xiommu1/oc8051_page_table_i/n611 , 
        \oc8051_xiommu1/oc8051_page_table_i/n612 , \oc8051_xiommu1/oc8051_page_table_i/n613 , 
        \oc8051_xiommu1/oc8051_page_table_i/n614 , \oc8051_xiommu1/oc8051_page_table_i/n615 , 
        \oc8051_xiommu1/oc8051_page_table_i/n616 , \oc8051_xiommu1/oc8051_page_table_i/n617 , 
        \oc8051_xiommu1/oc8051_page_table_i/n618 , \oc8051_xiommu1/oc8051_page_table_i/n619 , 
        \oc8051_xiommu1/oc8051_page_table_i/n620 , \oc8051_xiommu1/oc8051_page_table_i/n621 , 
        \oc8051_xiommu1/oc8051_page_table_i/n622 , \oc8051_xiommu1/oc8051_page_table_i/n623 , 
        \oc8051_xiommu1/oc8051_page_table_i/n624 , \oc8051_xiommu1/oc8051_page_table_i/n625 , 
        \oc8051_xiommu1/oc8051_page_table_i/n626 , \oc8051_xiommu1/oc8051_page_table_i/n627 , 
        \oc8051_xiommu1/oc8051_page_table_i/n628 , \oc8051_xiommu1/oc8051_page_table_i/n629 , 
        \oc8051_xiommu1/oc8051_page_table_i/n630 , \oc8051_xiommu1/oc8051_page_table_i/n631 , 
        \oc8051_xiommu1/oc8051_page_table_i/n632 , \oc8051_xiommu1/oc8051_page_table_i/n633 , 
        \oc8051_xiommu1/oc8051_page_table_i/n634 , \oc8051_xiommu1/oc8051_page_table_i/n635 , 
        \oc8051_xiommu1/oc8051_page_table_i/n636 , \oc8051_xiommu1/oc8051_page_table_i/n637 , 
        \oc8051_xiommu1/oc8051_page_table_i/n638 , \oc8051_xiommu1/oc8051_page_table_i/n639 , 
        \oc8051_xiommu1/oc8051_page_table_i/n640 , \oc8051_xiommu1/oc8051_page_table_i/n641 , 
        \oc8051_xiommu1/oc8051_page_table_i/n642 , \oc8051_xiommu1/oc8051_page_table_i/n643 , 
        \oc8051_xiommu1/oc8051_page_table_i/n644 , \oc8051_xiommu1/oc8051_page_table_i/n645 , 
        \oc8051_xiommu1/oc8051_page_table_i/n646 , \oc8051_xiommu1/oc8051_page_table_i/n647 , 
        \oc8051_xiommu1/oc8051_page_table_i/n648 , \oc8051_xiommu1/oc8051_page_table_i/n649 , 
        \oc8051_xiommu1/oc8051_page_table_i/n650 , \oc8051_xiommu1/oc8051_page_table_i/n651 , 
        \oc8051_xiommu1/oc8051_page_table_i/n652 , \oc8051_xiommu1/oc8051_page_table_i/n653 , 
        \oc8051_xiommu1/oc8051_page_table_i/n654 , \oc8051_xiommu1/oc8051_page_table_i/n655 , 
        \oc8051_xiommu1/oc8051_page_table_i/n656 , \oc8051_xiommu1/oc8051_page_table_i/n657 , 
        \oc8051_xiommu1/oc8051_page_table_i/n658 , \oc8051_xiommu1/oc8051_page_table_i/n659 , 
        \oc8051_xiommu1/oc8051_page_table_i/n660 , \oc8051_xiommu1/oc8051_page_table_i/n661 , 
        \oc8051_xiommu1/oc8051_page_table_i/n662 , \oc8051_xiommu1/oc8051_page_table_i/n663 , 
        \oc8051_xiommu1/oc8051_page_table_i/n664 , \oc8051_xiommu1/oc8051_page_table_i/n665 , 
        \oc8051_xiommu1/oc8051_page_table_i/n666 , \oc8051_xiommu1/oc8051_page_table_i/n667 , 
        \oc8051_xiommu1/oc8051_page_table_i/n668 , \oc8051_xiommu1/oc8051_page_table_i/n669 , 
        \oc8051_xiommu1/oc8051_page_table_i/n670 , \oc8051_xiommu1/oc8051_page_table_i/n671 , 
        \oc8051_xiommu1/oc8051_page_table_i/n672 , \oc8051_xiommu1/oc8051_page_table_i/n673 , 
        \oc8051_xiommu1/oc8051_page_table_i/n674 , \oc8051_xiommu1/oc8051_page_table_i/n675 , 
        \oc8051_xiommu1/oc8051_page_table_i/n676 , \oc8051_xiommu1/oc8051_page_table_i/n677 , 
        \oc8051_xiommu1/oc8051_page_table_i/n678 , \oc8051_xiommu1/oc8051_page_table_i/n679 , 
        \oc8051_xiommu1/oc8051_page_table_i/n680 , \oc8051_xiommu1/oc8051_page_table_i/n681 , 
        \oc8051_xiommu1/oc8051_page_table_i/n682 , \oc8051_xiommu1/oc8051_page_table_i/n683 , 
        \oc8051_xiommu1/oc8051_page_table_i/n684 , \oc8051_xiommu1/oc8051_page_table_i/n685 , 
        \oc8051_xiommu1/oc8051_page_table_i/n686 , \oc8051_xiommu1/oc8051_page_table_i/n687 , 
        \oc8051_xiommu1/oc8051_page_table_i/n688 , \oc8051_xiommu1/oc8051_page_table_i/n689 , 
        \oc8051_xiommu1/oc8051_page_table_i/n690 , \oc8051_xiommu1/oc8051_page_table_i/n691 , 
        \oc8051_xiommu1/oc8051_page_table_i/n692 , \oc8051_xiommu1/oc8051_page_table_i/n693 , 
        \oc8051_xiommu1/oc8051_page_table_i/n694 , \oc8051_xiommu1/oc8051_page_table_i/n695 , 
        \oc8051_xiommu1/oc8051_page_table_i/n696 , \oc8051_xiommu1/oc8051_page_table_i/n697 , 
        \oc8051_xiommu1/oc8051_page_table_i/n698 , \oc8051_xiommu1/oc8051_page_table_i/n699 , 
        \oc8051_xiommu1/oc8051_page_table_i/n700 , \oc8051_xiommu1/oc8051_page_table_i/n701 , 
        \oc8051_xiommu1/oc8051_page_table_i/n702 , \oc8051_xiommu1/oc8051_page_table_i/n703 , 
        \oc8051_xiommu1/oc8051_page_table_i/n704 , \oc8051_xiommu1/oc8051_page_table_i/n705 , 
        \oc8051_xiommu1/oc8051_page_table_i/n706 , \oc8051_xiommu1/oc8051_page_table_i/n707 , 
        \oc8051_xiommu1/oc8051_page_table_i/n708 , \oc8051_xiommu1/oc8051_page_table_i/n709 , 
        \oc8051_xiommu1/oc8051_page_table_i/n710 , \oc8051_xiommu1/oc8051_page_table_i/n711 , 
        \oc8051_xiommu1/oc8051_page_table_i/n712 , \oc8051_xiommu1/oc8051_page_table_i/n713 , 
        \oc8051_xiommu1/oc8051_page_table_i/n714 , \oc8051_xiommu1/oc8051_page_table_i/n715 , 
        \oc8051_xiommu1/oc8051_page_table_i/n716 , \oc8051_xiommu1/oc8051_page_table_i/n717 , 
        \oc8051_xiommu1/oc8051_page_table_i/n718 , \oc8051_xiommu1/oc8051_page_table_i/n719 , 
        \oc8051_xiommu1/oc8051_page_table_i/n720 , \oc8051_xiommu1/oc8051_page_table_i/n721 , 
        \oc8051_xiommu1/oc8051_page_table_i/n722 , \oc8051_xiommu1/oc8051_page_table_i/n723 , 
        \oc8051_xiommu1/oc8051_page_table_i/n724 , \oc8051_xiommu1/oc8051_page_table_i/n725 , 
        \oc8051_xiommu1/oc8051_page_table_i/n726 , \oc8051_xiommu1/oc8051_page_table_i/n727 , 
        \oc8051_xiommu1/oc8051_page_table_i/n728 , \oc8051_xiommu1/oc8051_page_table_i/n729 , 
        \oc8051_xiommu1/oc8051_page_table_i/n730 , \oc8051_xiommu1/oc8051_page_table_i/n731 , 
        \oc8051_xiommu1/oc8051_page_table_i/n732 , \oc8051_xiommu1/oc8051_page_table_i/n733 , 
        \oc8051_xiommu1/oc8051_page_table_i/n734 , \oc8051_xiommu1/oc8051_page_table_i/n735 , 
        \oc8051_xiommu1/oc8051_page_table_i/n736 , \oc8051_xiommu1/oc8051_page_table_i/n737 , 
        \oc8051_xiommu1/oc8051_page_table_i/n738 , \oc8051_xiommu1/oc8051_page_table_i/n739 , 
        \oc8051_xiommu1/oc8051_page_table_i/n740 , \oc8051_xiommu1/oc8051_page_table_i/n741 , 
        \oc8051_xiommu1/oc8051_page_table_i/n742 , \oc8051_xiommu1/oc8051_page_table_i/n743 , 
        \oc8051_xiommu1/oc8051_page_table_i/n744 , \oc8051_xiommu1/oc8051_page_table_i/n745 , 
        \oc8051_xiommu1/oc8051_page_table_i/n746 , \oc8051_xiommu1/oc8051_page_table_i/n747 , 
        \oc8051_xiommu1/oc8051_page_table_i/n748 , \oc8051_xiommu1/oc8051_page_table_i/n749 , 
        \oc8051_xiommu1/oc8051_page_table_i/n750 , \oc8051_xiommu1/oc8051_page_table_i/n751 , 
        \oc8051_xiommu1/oc8051_page_table_i/n752 , \oc8051_xiommu1/oc8051_page_table_i/n753 , 
        \oc8051_xiommu1/oc8051_page_table_i/n754 , \oc8051_xiommu1/oc8051_page_table_i/n755 , 
        \oc8051_xiommu1/oc8051_page_table_i/n756 , \oc8051_xiommu1/oc8051_page_table_i/n757 , 
        \oc8051_xiommu1/oc8051_page_table_i/n758 , \oc8051_xiommu1/oc8051_page_table_i/n759 , 
        \oc8051_xiommu1/oc8051_page_table_i/n760 , \oc8051_xiommu1/oc8051_page_table_i/n761 , 
        \oc8051_xiommu1/oc8051_page_table_i/n762 , \oc8051_xiommu1/oc8051_page_table_i/n763 , 
        \oc8051_xiommu1/oc8051_page_table_i/n764 , \oc8051_xiommu1/oc8051_page_table_i/n765 , 
        \oc8051_xiommu1/oc8051_page_table_i/n766 , \oc8051_xiommu1/oc8051_page_table_i/n767 , 
        \oc8051_xiommu1/oc8051_page_table_i/n768 , \oc8051_xiommu1/oc8051_page_table_i/n769 , 
        \oc8051_xiommu1/oc8051_page_table_i/n770 , \oc8051_xiommu1/oc8051_page_table_i/n771 , 
        \oc8051_xiommu1/oc8051_page_table_i/n772 , \oc8051_xiommu1/oc8051_page_table_i/n773 , 
        \oc8051_xiommu1/oc8051_page_table_i/n774 , \oc8051_xiommu1/oc8051_page_table_i/n775 , 
        \oc8051_xiommu1/oc8051_page_table_i/n776 , \oc8051_xiommu1/oc8051_page_table_i/n777 , 
        \oc8051_xiommu1/oc8051_page_table_i/n778 , \oc8051_xiommu1/oc8051_page_table_i/n779 , 
        \oc8051_xiommu1/oc8051_page_table_i/n780 , \oc8051_xiommu1/oc8051_page_table_i/n781 , 
        \oc8051_xiommu1/oc8051_page_table_i/n782 , \oc8051_xiommu1/oc8051_page_table_i/n783 , 
        \oc8051_xiommu1/oc8051_page_table_i/n784 , \oc8051_xiommu1/oc8051_page_table_i/n785 , 
        \oc8051_xiommu1/oc8051_page_table_i/n786 , \oc8051_xiommu1/oc8051_page_table_i/n787 , 
        \oc8051_xiommu1/oc8051_page_table_i/n788 , \oc8051_xiommu1/oc8051_page_table_i/n789 , 
        \oc8051_xiommu1/oc8051_page_table_i/n790 , \oc8051_xiommu1/oc8051_page_table_i/n791 , 
        \oc8051_xiommu1/oc8051_page_table_i/n792 , \oc8051_xiommu1/oc8051_page_table_i/n793 , 
        \oc8051_xiommu1/oc8051_page_table_i/n794 , \oc8051_xiommu1/oc8051_page_table_i/n795 , 
        \oc8051_xiommu1/oc8051_page_table_i/n796 , \oc8051_xiommu1/oc8051_page_table_i/n797 , 
        \oc8051_xiommu1/oc8051_page_table_i/n798 , \oc8051_xiommu1/oc8051_page_table_i/n799 , 
        \oc8051_xiommu1/oc8051_page_table_i/n800 , \oc8051_xiommu1/oc8051_page_table_i/n801 , 
        \oc8051_xiommu1/oc8051_page_table_i/n802 , \oc8051_xiommu1/oc8051_page_table_i/n803 , 
        \oc8051_xiommu1/oc8051_page_table_i/n804 , \oc8051_xiommu1/oc8051_page_table_i/n805 , 
        \oc8051_xiommu1/oc8051_page_table_i/n806 , \oc8051_xiommu1/oc8051_page_table_i/n807 , 
        \oc8051_xiommu1/oc8051_page_table_i/n808 , \oc8051_xiommu1/oc8051_page_table_i/n809 , 
        \oc8051_xiommu1/oc8051_page_table_i/n810 , \oc8051_xiommu1/oc8051_page_table_i/n811 , 
        \oc8051_xiommu1/oc8051_page_table_i/n812 , \oc8051_xiommu1/oc8051_page_table_i/n813 , 
        \oc8051_xiommu1/oc8051_page_table_i/n814 , \oc8051_xiommu1/oc8051_page_table_i/n815 , 
        \oc8051_xiommu1/oc8051_page_table_i/n816 , \oc8051_xiommu1/oc8051_page_table_i/n817 , 
        \oc8051_xiommu1/oc8051_page_table_i/n818 , \oc8051_xiommu1/oc8051_page_table_i/n819 , 
        \oc8051_xiommu1/oc8051_page_table_i/n820 , \oc8051_xiommu1/oc8051_page_table_i/n821 , 
        \oc8051_xiommu1/oc8051_page_table_i/n822 , \oc8051_xiommu1/oc8051_page_table_i/n823 , 
        \oc8051_xiommu1/oc8051_page_table_i/n824 , \oc8051_xiommu1/oc8051_page_table_i/n825 , 
        \oc8051_xiommu1/oc8051_page_table_i/n826 , \oc8051_xiommu1/oc8051_page_table_i/n827 , 
        \oc8051_xiommu1/oc8051_page_table_i/n828 , \oc8051_xiommu1/oc8051_page_table_i/n829 , 
        \oc8051_xiommu1/oc8051_page_table_i/n830 , \oc8051_xiommu1/oc8051_page_table_i/n831 , 
        \oc8051_xiommu1/oc8051_page_table_i/n832 , \oc8051_xiommu1/oc8051_page_table_i/n833 , 
        \oc8051_xiommu1/oc8051_page_table_i/n834 , \oc8051_xiommu1/oc8051_page_table_i/n835 , 
        \oc8051_xiommu1/oc8051_page_table_i/n836 , \oc8051_xiommu1/oc8051_page_table_i/n837 , 
        \oc8051_xiommu1/oc8051_page_table_i/n838 , \oc8051_xiommu1/oc8051_page_table_i/n839 , 
        \oc8051_xiommu1/oc8051_page_table_i/n840 , \oc8051_xiommu1/oc8051_page_table_i/n841 , 
        \oc8051_xiommu1/oc8051_page_table_i/n842 , \oc8051_xiommu1/oc8051_page_table_i/n843 , 
        \oc8051_xiommu1/oc8051_page_table_i/n844 , \oc8051_xiommu1/oc8051_page_table_i/n845 , 
        \oc8051_xiommu1/oc8051_page_table_i/n846 , \oc8051_xiommu1/oc8051_page_table_i/n847 , 
        \oc8051_xiommu1/oc8051_page_table_i/n848 , \oc8051_xiommu1/oc8051_page_table_i/n849 , 
        \oc8051_xiommu1/oc8051_page_table_i/n850 , \oc8051_xiommu1/oc8051_page_table_i/n851 , 
        \oc8051_xiommu1/oc8051_page_table_i/n852 , \oc8051_xiommu1/oc8051_page_table_i/n853 , 
        \oc8051_xiommu1/oc8051_page_table_i/n854 , \oc8051_xiommu1/oc8051_page_table_i/n855 , 
        \oc8051_xiommu1/oc8051_page_table_i/n856 , \oc8051_xiommu1/oc8051_page_table_i/n857 , 
        \oc8051_xiommu1/oc8051_page_table_i/n858 , \oc8051_xiommu1/oc8051_page_table_i/n859 , 
        \oc8051_xiommu1/oc8051_page_table_i/n860 , \oc8051_xiommu1/oc8051_page_table_i/n861 , 
        \oc8051_xiommu1/oc8051_page_table_i/n862 , \oc8051_xiommu1/oc8051_page_table_i/n863 , 
        \oc8051_xiommu1/oc8051_page_table_i/n864 , \oc8051_xiommu1/oc8051_page_table_i/n865 , 
        \oc8051_xiommu1/oc8051_page_table_i/n866 , \oc8051_xiommu1/oc8051_page_table_i/n867 , 
        \oc8051_xiommu1/oc8051_page_table_i/n868 , \oc8051_xiommu1/oc8051_page_table_i/n869 , 
        \oc8051_xiommu1/oc8051_page_table_i/n870 , \oc8051_xiommu1/oc8051_page_table_i/n871 , 
        \oc8051_xiommu1/oc8051_page_table_i/n872 , \oc8051_xiommu1/oc8051_page_table_i/n873 , 
        \oc8051_xiommu1/oc8051_page_table_i/n874 , \oc8051_xiommu1/oc8051_page_table_i/n875 , 
        \oc8051_xiommu1/oc8051_page_table_i/n876 , \oc8051_xiommu1/oc8051_page_table_i/n877 , 
        \oc8051_xiommu1/oc8051_page_table_i/n878 , \oc8051_xiommu1/oc8051_page_table_i/n879 , 
        \oc8051_xiommu1/oc8051_page_table_i/n880 , \oc8051_xiommu1/oc8051_page_table_i/n881 , 
        \oc8051_xiommu1/oc8051_page_table_i/n882 , \oc8051_xiommu1/oc8051_page_table_i/n883 , 
        \oc8051_xiommu1/oc8051_page_table_i/n884 , \oc8051_xiommu1/oc8051_page_table_i/n885 , 
        \oc8051_xiommu1/oc8051_page_table_i/n886 , \oc8051_xiommu1/oc8051_page_table_i/n887 , 
        \oc8051_xiommu1/oc8051_page_table_i/n888 , \oc8051_xiommu1/oc8051_page_table_i/n889 , 
        \oc8051_xiommu1/oc8051_page_table_i/n890 , \oc8051_xiommu1/oc8051_page_table_i/n891 , 
        \oc8051_xiommu1/oc8051_page_table_i/n892 , \oc8051_xiommu1/oc8051_page_table_i/n893 , 
        \oc8051_xiommu1/oc8051_page_table_i/n894 , \oc8051_xiommu1/oc8051_page_table_i/n895 , 
        \oc8051_xiommu1/oc8051_page_table_i/n896 , \oc8051_xiommu1/oc8051_page_table_i/n897 , 
        \oc8051_xiommu1/oc8051_page_table_i/n898 , \oc8051_xiommu1/oc8051_page_table_i/n899 , 
        \oc8051_xiommu1/oc8051_page_table_i/n900 , \oc8051_xiommu1/oc8051_page_table_i/n901 , 
        \oc8051_xiommu1/oc8051_page_table_i/n902 , \oc8051_xiommu1/oc8051_page_table_i/n903 , 
        \oc8051_xiommu1/oc8051_page_table_i/n904 , \oc8051_xiommu1/oc8051_page_table_i/n905 , 
        \oc8051_xiommu1/oc8051_page_table_i/n906 , \oc8051_xiommu1/oc8051_page_table_i/n907 , 
        \oc8051_xiommu1/oc8051_page_table_i/n908 , \oc8051_xiommu1/oc8051_page_table_i/n909 , 
        \oc8051_xiommu1/oc8051_page_table_i/n910 , \oc8051_xiommu1/oc8051_page_table_i/n911 , 
        \oc8051_xiommu1/oc8051_page_table_i/n912 , \oc8051_xiommu1/oc8051_page_table_i/n913 , 
        \oc8051_xiommu1/oc8051_page_table_i/n914 , \oc8051_xiommu1/oc8051_page_table_i/n915 , 
        \oc8051_xiommu1/oc8051_page_table_i/n916 , \oc8051_xiommu1/oc8051_page_table_i/n917 , 
        \oc8051_xiommu1/oc8051_page_table_i/n918 , \oc8051_xiommu1/oc8051_page_table_i/n919 , 
        \oc8051_xiommu1/oc8051_page_table_i/n920 , \oc8051_xiommu1/oc8051_page_table_i/n921 , 
        \oc8051_xiommu1/oc8051_page_table_i/n922 , \oc8051_xiommu1/oc8051_page_table_i/n923 , 
        \oc8051_xiommu1/oc8051_page_table_i/n924 , \oc8051_xiommu1/oc8051_page_table_i/n925 , 
        \oc8051_xiommu1/oc8051_page_table_i/n926 , \oc8051_xiommu1/oc8051_page_table_i/n927 , 
        \oc8051_xiommu1/oc8051_page_table_i/n928 , \oc8051_xiommu1/oc8051_page_table_i/n929 , 
        \oc8051_xiommu1/oc8051_page_table_i/n930 , \oc8051_xiommu1/oc8051_page_table_i/n931 , 
        \oc8051_xiommu1/oc8051_page_table_i/n932 , \oc8051_xiommu1/oc8051_page_table_i/n933 , 
        \oc8051_xiommu1/oc8051_page_table_i/n934 , \oc8051_xiommu1/oc8051_page_table_i/n935 , 
        \oc8051_xiommu1/oc8051_page_table_i/n936 , \oc8051_xiommu1/oc8051_page_table_i/n937 , 
        \oc8051_xiommu1/oc8051_page_table_i/n938 , \oc8051_xiommu1/oc8051_page_table_i/n939 , 
        \oc8051_xiommu1/oc8051_page_table_i/n940 , \oc8051_xiommu1/oc8051_page_table_i/n941 , 
        \oc8051_xiommu1/oc8051_page_table_i/n942 , \oc8051_xiommu1/oc8051_page_table_i/n943 , 
        \oc8051_xiommu1/oc8051_page_table_i/n944 , \oc8051_xiommu1/oc8051_page_table_i/n945 , 
        \oc8051_xiommu1/oc8051_page_table_i/n946 , \oc8051_xiommu1/oc8051_page_table_i/n947 , 
        \oc8051_xiommu1/oc8051_page_table_i/n948 , \oc8051_xiommu1/oc8051_page_table_i/n949 , 
        \oc8051_xiommu1/oc8051_page_table_i/n950 , \oc8051_xiommu1/oc8051_page_table_i/n951 , 
        \oc8051_xiommu1/oc8051_page_table_i/n952 , \oc8051_xiommu1/oc8051_page_table_i/n953 , 
        \oc8051_xiommu1/oc8051_page_table_i/n954 , \oc8051_xiommu1/oc8051_page_table_i/n955 , 
        \oc8051_xiommu1/oc8051_page_table_i/n956 , \oc8051_xiommu1/oc8051_page_table_i/n957 , 
        \oc8051_xiommu1/oc8051_page_table_i/n958 , \oc8051_xiommu1/oc8051_page_table_i/n959 , 
        \oc8051_xiommu1/oc8051_page_table_i/n960 , \oc8051_xiommu1/oc8051_page_table_i/n961 , 
        \oc8051_xiommu1/oc8051_page_table_i/n962 , \oc8051_xiommu1/oc8051_page_table_i/n963 , 
        \oc8051_xiommu1/oc8051_page_table_i/n964 , \oc8051_xiommu1/oc8051_page_table_i/n965 , 
        \oc8051_xiommu1/oc8051_page_table_i/n966 , \oc8051_xiommu1/oc8051_page_table_i/n967 , 
        \oc8051_xiommu1/oc8051_page_table_i/n968 , \oc8051_xiommu1/oc8051_page_table_i/n969 , 
        \oc8051_xiommu1/oc8051_page_table_i/n970 , \oc8051_xiommu1/oc8051_page_table_i/n971 , 
        \oc8051_xiommu1/oc8051_page_table_i/n972 , \oc8051_xiommu1/oc8051_page_table_i/n973 , 
        \oc8051_xiommu1/oc8051_page_table_i/n974 , \oc8051_xiommu1/oc8051_page_table_i/n975 , 
        \oc8051_xiommu1/oc8051_page_table_i/n976 , \oc8051_xiommu1/oc8051_page_table_i/n977 , 
        \oc8051_xiommu1/oc8051_page_table_i/n978 , \oc8051_xiommu1/oc8051_page_table_i/n979 , 
        \oc8051_xiommu1/oc8051_page_table_i/n980 , \oc8051_xiommu1/oc8051_page_table_i/n981 , 
        \oc8051_xiommu1/oc8051_page_table_i/n982 , \oc8051_xiommu1/oc8051_page_table_i/n983 , 
        \oc8051_xiommu1/oc8051_page_table_i/n984 , \oc8051_xiommu1/oc8051_page_table_i/n985 , 
        \oc8051_xiommu1/oc8051_page_table_i/n986 , \oc8051_xiommu1/oc8051_page_table_i/n987 , 
        \oc8051_xiommu1/oc8051_page_table_i/n988 , \oc8051_xiommu1/oc8051_page_table_i/n989 , 
        \oc8051_xiommu1/oc8051_page_table_i/n990 , \oc8051_xiommu1/oc8051_page_table_i/n991 , 
        \oc8051_xiommu1/oc8051_page_table_i/n992 , \oc8051_xiommu1/oc8051_page_table_i/n993 , 
        \oc8051_xiommu1/oc8051_page_table_i/n994 , \oc8051_xiommu1/oc8051_page_table_i/n995 , 
        \oc8051_xiommu1/oc8051_page_table_i/n996 , \oc8051_xiommu1/oc8051_page_table_i/n997 , 
        \oc8051_xiommu1/oc8051_page_table_i/n998 , \oc8051_xiommu1/oc8051_page_table_i/n999 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1000 , \oc8051_xiommu1/oc8051_page_table_i/n1001 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1002 , \oc8051_xiommu1/oc8051_page_table_i/n1003 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1004 , \oc8051_xiommu1/oc8051_page_table_i/n1005 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1006 , \oc8051_xiommu1/oc8051_page_table_i/n1007 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1008 , \oc8051_xiommu1/oc8051_page_table_i/n1009 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1010 , \oc8051_xiommu1/oc8051_page_table_i/n1011 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1012 , \oc8051_xiommu1/oc8051_page_table_i/n1013 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1014 , \oc8051_xiommu1/oc8051_page_table_i/n1015 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1016 , \oc8051_xiommu1/oc8051_page_table_i/n1017 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1018 , \oc8051_xiommu1/oc8051_page_table_i/n1019 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1020 , \oc8051_xiommu1/oc8051_page_table_i/n1021 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1022 , \oc8051_xiommu1/oc8051_page_table_i/n1023 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1024 , \oc8051_xiommu1/oc8051_page_table_i/n1025 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1026 , \oc8051_xiommu1/oc8051_page_table_i/n1027 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1028 , \oc8051_xiommu1/oc8051_page_table_i/n1029 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1030 , \oc8051_xiommu1/oc8051_page_table_i/n1031 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1032 , \oc8051_xiommu1/oc8051_page_table_i/n1033 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1034 , \oc8051_xiommu1/oc8051_page_table_i/n1035 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1036 , \oc8051_xiommu1/oc8051_page_table_i/n1037 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1038 , \oc8051_xiommu1/oc8051_page_table_i/n1039 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1040 , \oc8051_xiommu1/oc8051_page_table_i/n1041 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1042 , \oc8051_xiommu1/oc8051_page_table_i/n1043 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1044 , \oc8051_xiommu1/oc8051_page_table_i/n1045 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1046 , \oc8051_xiommu1/oc8051_page_table_i/n1047 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1048 , \oc8051_xiommu1/oc8051_page_table_i/n1049 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1050 , \oc8051_xiommu1/oc8051_page_table_i/n1051 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1052 , \oc8051_xiommu1/oc8051_page_table_i/n1053 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1054 , \oc8051_xiommu1/oc8051_page_table_i/n1055 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1056 , \oc8051_xiommu1/oc8051_page_table_i/n1057 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1058 , \oc8051_xiommu1/oc8051_page_table_i/n1059 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1060 , \oc8051_xiommu1/oc8051_page_table_i/n1061 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1062 , \oc8051_xiommu1/oc8051_page_table_i/n1063 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1064 , \oc8051_xiommu1/oc8051_page_table_i/n1065 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1066 , \oc8051_xiommu1/oc8051_page_table_i/n1067 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1068 , \oc8051_xiommu1/oc8051_page_table_i/n1069 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1070 , \oc8051_xiommu1/oc8051_page_table_i/n1071 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1072 , \oc8051_xiommu1/oc8051_page_table_i/n1073 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1074 , \oc8051_xiommu1/oc8051_page_table_i/n1075 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1076 , \oc8051_xiommu1/oc8051_page_table_i/n1077 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1078 , \oc8051_xiommu1/oc8051_page_table_i/n1079 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1080 , \oc8051_xiommu1/oc8051_page_table_i/n1081 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1082 , \oc8051_xiommu1/oc8051_page_table_i/n1083 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1084 , \oc8051_xiommu1/oc8051_page_table_i/n1085 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1086 , \oc8051_xiommu1/oc8051_page_table_i/n1087 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1088 , \oc8051_xiommu1/oc8051_page_table_i/n1089 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1090 , \oc8051_xiommu1/oc8051_page_table_i/n1091 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1092 , \oc8051_xiommu1/oc8051_page_table_i/n1093 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1094 , \oc8051_xiommu1/oc8051_page_table_i/n1095 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1096 , \oc8051_xiommu1/oc8051_page_table_i/n1097 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1098 , \oc8051_xiommu1/oc8051_page_table_i/n1099 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1100 , \oc8051_xiommu1/oc8051_page_table_i/n1101 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1102 , \oc8051_xiommu1/oc8051_page_table_i/n1103 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1104 , \oc8051_xiommu1/oc8051_page_table_i/n1105 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1106 , \oc8051_xiommu1/oc8051_page_table_i/n1107 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1108 , \oc8051_xiommu1/oc8051_page_table_i/n1109 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1110 , \oc8051_xiommu1/oc8051_page_table_i/n1111 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1112 , \oc8051_xiommu1/oc8051_page_table_i/n1113 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1114 , \oc8051_xiommu1/oc8051_page_table_i/n1115 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1116 , \oc8051_xiommu1/oc8051_page_table_i/n1117 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1118 , \oc8051_xiommu1/oc8051_page_table_i/n1119 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1120 , \oc8051_xiommu1/oc8051_page_table_i/n1121 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1122 , \oc8051_xiommu1/oc8051_page_table_i/n1123 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1124 , \oc8051_xiommu1/oc8051_page_table_i/n1125 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1126 , \oc8051_xiommu1/oc8051_page_table_i/n1127 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1128 , \oc8051_xiommu1/oc8051_page_table_i/n1129 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1130 , \oc8051_xiommu1/oc8051_page_table_i/n1131 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1132 , \oc8051_xiommu1/oc8051_page_table_i/n1133 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1134 , \oc8051_xiommu1/oc8051_page_table_i/n1135 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1136 , \oc8051_xiommu1/oc8051_page_table_i/n1137 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1138 , \oc8051_xiommu1/oc8051_page_table_i/n1139 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1140 , \oc8051_xiommu1/oc8051_page_table_i/n1141 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1142 , \oc8051_xiommu1/oc8051_page_table_i/n1143 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1144 , \oc8051_xiommu1/oc8051_page_table_i/n1145 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1146 , \oc8051_xiommu1/oc8051_page_table_i/n1147 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1148 , \oc8051_xiommu1/oc8051_page_table_i/n1149 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1150 , \oc8051_xiommu1/oc8051_page_table_i/n1151 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1152 , \oc8051_xiommu1/oc8051_page_table_i/n1153 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1154 , \oc8051_xiommu1/oc8051_page_table_i/n1155 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1156 , \oc8051_xiommu1/oc8051_page_table_i/n1157 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1158 , \oc8051_xiommu1/oc8051_page_table_i/n1159 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1160 , \oc8051_xiommu1/oc8051_page_table_i/n1161 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1162 , \oc8051_xiommu1/oc8051_page_table_i/n1163 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1164 , \oc8051_xiommu1/oc8051_page_table_i/n1165 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1166 , \oc8051_xiommu1/oc8051_page_table_i/n1167 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1168 , \oc8051_xiommu1/oc8051_page_table_i/n1169 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1170 , \oc8051_xiommu1/oc8051_page_table_i/n1171 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1172 , \oc8051_xiommu1/oc8051_page_table_i/n1173 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1174 , \oc8051_xiommu1/oc8051_page_table_i/n1175 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1176 , \oc8051_xiommu1/oc8051_page_table_i/n1177 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1178 , \oc8051_xiommu1/oc8051_page_table_i/n1179 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1180 , \oc8051_xiommu1/oc8051_page_table_i/n1181 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1182 , \oc8051_xiommu1/oc8051_page_table_i/n1183 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1184 , \oc8051_xiommu1/oc8051_page_table_i/n1185 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1186 , \oc8051_xiommu1/oc8051_page_table_i/n1187 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1188 , \oc8051_xiommu1/oc8051_page_table_i/n1189 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1190 , \oc8051_xiommu1/oc8051_page_table_i/n1191 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1192 , \oc8051_xiommu1/oc8051_page_table_i/n1193 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1194 , \oc8051_xiommu1/oc8051_page_table_i/n1195 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1196 , \oc8051_xiommu1/oc8051_page_table_i/n1197 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1198 , \oc8051_xiommu1/oc8051_page_table_i/n1199 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1200 , \oc8051_xiommu1/oc8051_page_table_i/n1201 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1202 , \oc8051_xiommu1/oc8051_page_table_i/n1203 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1204 , \oc8051_xiommu1/oc8051_page_table_i/n1205 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1206 , \oc8051_xiommu1/oc8051_page_table_i/n1207 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1208 , \oc8051_xiommu1/oc8051_page_table_i/n1209 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1210 , \oc8051_xiommu1/oc8051_page_table_i/n1211 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1212 , \oc8051_xiommu1/oc8051_page_table_i/n1213 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1214 , \oc8051_xiommu1/oc8051_page_table_i/n1215 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1216 , \oc8051_xiommu1/oc8051_page_table_i/n1217 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1218 , \oc8051_xiommu1/oc8051_page_table_i/n1219 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1220 , \oc8051_xiommu1/oc8051_page_table_i/n1221 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1222 , \oc8051_xiommu1/oc8051_page_table_i/n1223 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1224 , \oc8051_xiommu1/oc8051_page_table_i/n1225 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1226 , \oc8051_xiommu1/oc8051_page_table_i/n1227 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1228 , \oc8051_xiommu1/oc8051_page_table_i/n1229 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1230 , \oc8051_xiommu1/oc8051_page_table_i/n1231 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1232 , \oc8051_xiommu1/oc8051_page_table_i/n1233 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1234 , \oc8051_xiommu1/oc8051_page_table_i/n1235 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1236 , \oc8051_xiommu1/oc8051_page_table_i/n1237 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1238 , \oc8051_xiommu1/oc8051_page_table_i/n1239 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1240 , \oc8051_xiommu1/oc8051_page_table_i/n1241 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1242 , \oc8051_xiommu1/oc8051_page_table_i/n1243 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1244 , \oc8051_xiommu1/oc8051_page_table_i/n1245 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1246 , \oc8051_xiommu1/oc8051_page_table_i/n1247 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1248 , \oc8051_xiommu1/oc8051_page_table_i/n1249 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1250 , \oc8051_xiommu1/oc8051_page_table_i/n1251 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1252 , \oc8051_xiommu1/oc8051_page_table_i/n1253 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1254 , \oc8051_xiommu1/oc8051_page_table_i/n1255 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1256 , \oc8051_xiommu1/oc8051_page_table_i/n1257 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1258 , \oc8051_xiommu1/oc8051_page_table_i/n1259 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1260 , \oc8051_xiommu1/oc8051_page_table_i/n1261 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1262 , \oc8051_xiommu1/oc8051_page_table_i/n1263 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1264 , \oc8051_xiommu1/oc8051_page_table_i/n1265 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1266 , \oc8051_xiommu1/oc8051_page_table_i/n1267 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1268 , \oc8051_xiommu1/oc8051_page_table_i/n1269 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1270 , \oc8051_xiommu1/oc8051_page_table_i/n1271 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1272 , \oc8051_xiommu1/oc8051_page_table_i/n1273 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1274 , \oc8051_xiommu1/oc8051_page_table_i/n1275 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1276 , \oc8051_xiommu1/oc8051_page_table_i/n1277 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1278 , \oc8051_xiommu1/oc8051_page_table_i/n1279 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1280 , \oc8051_xiommu1/oc8051_page_table_i/n1281 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1282 , \oc8051_xiommu1/oc8051_page_table_i/n1283 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1284 , \oc8051_xiommu1/oc8051_page_table_i/n1285 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1286 , \oc8051_xiommu1/oc8051_page_table_i/n1287 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1288 , \oc8051_xiommu1/oc8051_page_table_i/n1289 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1290 , \oc8051_xiommu1/oc8051_page_table_i/n1291 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1292 , \oc8051_xiommu1/oc8051_page_table_i/n1293 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1294 , \oc8051_xiommu1/oc8051_page_table_i/n1295 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1296 , \oc8051_xiommu1/oc8051_page_table_i/n1297 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1298 , \oc8051_xiommu1/oc8051_page_table_i/n1299 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1300 , \oc8051_xiommu1/oc8051_page_table_i/n1301 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1302 , \oc8051_xiommu1/oc8051_page_table_i/n1303 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1304 , \oc8051_xiommu1/oc8051_page_table_i/n1305 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1306 , \oc8051_xiommu1/oc8051_page_table_i/n1307 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1308 , \oc8051_xiommu1/oc8051_page_table_i/n1309 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1310 , \oc8051_xiommu1/oc8051_page_table_i/n1311 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1312 , \oc8051_xiommu1/oc8051_page_table_i/n1313 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1314 , \oc8051_xiommu1/oc8051_page_table_i/n1315 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1316 , \oc8051_xiommu1/oc8051_page_table_i/n1317 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1318 , \oc8051_xiommu1/oc8051_page_table_i/n1319 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1320 , \oc8051_xiommu1/oc8051_page_table_i/n1321 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1322 , \oc8051_xiommu1/oc8051_page_table_i/n1323 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1324 , \oc8051_xiommu1/oc8051_page_table_i/n1325 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1326 , \oc8051_xiommu1/oc8051_page_table_i/n1327 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1328 , \oc8051_xiommu1/oc8051_page_table_i/n1329 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1330 , \oc8051_xiommu1/oc8051_page_table_i/n1331 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1332 , \oc8051_xiommu1/oc8051_page_table_i/n1333 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1334 , \oc8051_xiommu1/oc8051_page_table_i/n1335 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1336 , \oc8051_xiommu1/oc8051_page_table_i/n1337 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1338 , \oc8051_xiommu1/oc8051_page_table_i/n1339 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1340 , \oc8051_xiommu1/oc8051_page_table_i/n1341 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1342 , \oc8051_xiommu1/oc8051_page_table_i/n1343 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1344 , \oc8051_xiommu1/oc8051_page_table_i/n1345 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1346 , \oc8051_xiommu1/oc8051_page_table_i/n1347 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1348 , \oc8051_xiommu1/oc8051_page_table_i/n1349 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1350 , \oc8051_xiommu1/oc8051_page_table_i/n1351 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1352 , \oc8051_xiommu1/oc8051_page_table_i/n1353 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1354 , \oc8051_xiommu1/oc8051_page_table_i/n1355 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1356 , \oc8051_xiommu1/oc8051_page_table_i/n1357 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1358 , \oc8051_xiommu1/oc8051_page_table_i/n1359 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1360 , \oc8051_xiommu1/oc8051_page_table_i/n1361 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1362 , \oc8051_xiommu1/oc8051_page_table_i/n1363 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1364 , \oc8051_xiommu1/oc8051_page_table_i/n1365 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1366 , \oc8051_xiommu1/oc8051_page_table_i/n1367 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1368 , \oc8051_xiommu1/oc8051_page_table_i/n1369 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1370 , \oc8051_xiommu1/oc8051_page_table_i/n1371 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1372 , \oc8051_xiommu1/oc8051_page_table_i/n1373 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1374 , \oc8051_xiommu1/oc8051_page_table_i/n1375 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1376 , \oc8051_xiommu1/oc8051_page_table_i/n1377 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1378 , \oc8051_xiommu1/oc8051_page_table_i/n1379 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1380 , \oc8051_xiommu1/oc8051_page_table_i/n1381 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1382 , \oc8051_xiommu1/oc8051_page_table_i/n1383 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1384 , \oc8051_xiommu1/oc8051_page_table_i/n1385 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1386 , \oc8051_xiommu1/oc8051_page_table_i/n1387 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1388 , \oc8051_xiommu1/oc8051_page_table_i/n1389 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1390 , \oc8051_xiommu1/oc8051_page_table_i/n1391 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1392 , \oc8051_xiommu1/oc8051_page_table_i/n1393 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1394 , \oc8051_xiommu1/oc8051_page_table_i/n1395 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1396 , \oc8051_xiommu1/oc8051_page_table_i/n1397 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1398 , \oc8051_xiommu1/oc8051_page_table_i/n1399 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1400 , \oc8051_xiommu1/oc8051_page_table_i/n1401 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1402 , \oc8051_xiommu1/oc8051_page_table_i/n1403 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1404 , \oc8051_xiommu1/oc8051_page_table_i/n1405 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1406 , \oc8051_xiommu1/oc8051_page_table_i/n1407 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1408 , \oc8051_xiommu1/oc8051_page_table_i/n1409 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1410 , \oc8051_xiommu1/oc8051_page_table_i/n1411 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1412 , \oc8051_xiommu1/oc8051_page_table_i/n1413 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1414 , \oc8051_xiommu1/oc8051_page_table_i/n1415 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1416 , \oc8051_xiommu1/oc8051_page_table_i/n1417 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1418 , \oc8051_xiommu1/oc8051_page_table_i/n1419 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1420 , \oc8051_xiommu1/oc8051_page_table_i/n1421 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1422 , \oc8051_xiommu1/oc8051_page_table_i/n1423 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1424 , \oc8051_xiommu1/oc8051_page_table_i/n1425 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1426 , \oc8051_xiommu1/oc8051_page_table_i/n1427 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1428 , \oc8051_xiommu1/oc8051_page_table_i/n1429 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1430 , \oc8051_xiommu1/oc8051_page_table_i/n1431 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1432 , \oc8051_xiommu1/oc8051_page_table_i/n1433 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1434 , \oc8051_xiommu1/oc8051_page_table_i/n1435 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1436 , \oc8051_xiommu1/oc8051_page_table_i/n1437 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1438 , \oc8051_xiommu1/oc8051_page_table_i/n1439 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1440 , \oc8051_xiommu1/oc8051_page_table_i/n1441 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1442 , \oc8051_xiommu1/oc8051_page_table_i/n1443 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1444 , \oc8051_xiommu1/oc8051_page_table_i/n1445 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1446 , \oc8051_xiommu1/oc8051_page_table_i/n1447 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1448 , \oc8051_xiommu1/oc8051_page_table_i/n1449 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1450 , \oc8051_xiommu1/oc8051_page_table_i/n1451 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1452 , \oc8051_xiommu1/oc8051_page_table_i/n1453 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1454 , \oc8051_xiommu1/oc8051_page_table_i/n1455 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1456 , \oc8051_xiommu1/oc8051_page_table_i/n1457 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1458 , \oc8051_xiommu1/oc8051_page_table_i/n1459 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1460 , \oc8051_xiommu1/oc8051_page_table_i/n1461 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1462 , \oc8051_xiommu1/oc8051_page_table_i/n1463 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1464 , \oc8051_xiommu1/oc8051_page_table_i/n1465 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1466 , \oc8051_xiommu1/oc8051_page_table_i/n1467 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1468 , \oc8051_xiommu1/oc8051_page_table_i/n1469 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1470 , \oc8051_xiommu1/oc8051_page_table_i/n1471 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1472 , \oc8051_xiommu1/oc8051_page_table_i/n1473 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1474 , \oc8051_xiommu1/oc8051_page_table_i/n1475 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1476 , \oc8051_xiommu1/oc8051_page_table_i/n1477 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1478 , \oc8051_xiommu1/oc8051_page_table_i/n1479 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1480 , \oc8051_xiommu1/oc8051_page_table_i/n1481 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1482 , \oc8051_xiommu1/oc8051_page_table_i/n1483 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1484 , \oc8051_xiommu1/oc8051_page_table_i/n1485 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1486 , \oc8051_xiommu1/oc8051_page_table_i/n1487 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1488 , \oc8051_xiommu1/oc8051_page_table_i/n1489 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1490 , \oc8051_xiommu1/oc8051_page_table_i/n1491 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1492 , \oc8051_xiommu1/oc8051_page_table_i/n1493 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1494 , \oc8051_xiommu1/oc8051_page_table_i/n1495 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1496 , \oc8051_xiommu1/oc8051_page_table_i/n1497 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1498 , \oc8051_xiommu1/oc8051_page_table_i/n1499 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1500 , \oc8051_xiommu1/oc8051_page_table_i/n1501 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1502 , \oc8051_xiommu1/oc8051_page_table_i/n1503 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1504 , \oc8051_xiommu1/oc8051_page_table_i/n1505 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1506 , \oc8051_xiommu1/oc8051_page_table_i/n1507 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1508 , \oc8051_xiommu1/oc8051_page_table_i/n1509 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1510 , \oc8051_xiommu1/oc8051_page_table_i/n1511 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1512 , \oc8051_xiommu1/oc8051_page_table_i/n1513 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1514 , \oc8051_xiommu1/oc8051_page_table_i/n1515 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1516 , \oc8051_xiommu1/oc8051_page_table_i/n1517 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1518 , \oc8051_xiommu1/oc8051_page_table_i/n1519 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1520 , \oc8051_xiommu1/oc8051_page_table_i/n1521 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1522 , \oc8051_xiommu1/oc8051_page_table_i/n1523 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1524 , \oc8051_xiommu1/oc8051_page_table_i/n1525 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1526 , \oc8051_xiommu1/oc8051_page_table_i/n1527 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1528 , \oc8051_xiommu1/oc8051_page_table_i/n1529 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1530 , \oc8051_xiommu1/oc8051_page_table_i/n1531 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1532 , \oc8051_xiommu1/oc8051_page_table_i/n1533 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1534 , \oc8051_xiommu1/oc8051_page_table_i/n1535 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1536 , \oc8051_xiommu1/oc8051_page_table_i/n1537 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1538 , \oc8051_xiommu1/oc8051_page_table_i/n1539 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1540 , \oc8051_xiommu1/oc8051_page_table_i/n1541 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1542 , \oc8051_xiommu1/oc8051_page_table_i/n1543 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1544 , \oc8051_xiommu1/oc8051_page_table_i/n1545 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1546 , \oc8051_xiommu1/oc8051_page_table_i/n1547 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1548 , \oc8051_xiommu1/oc8051_page_table_i/n1549 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1550 , \oc8051_xiommu1/oc8051_page_table_i/n1551 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1552 , \oc8051_xiommu1/oc8051_page_table_i/n1553 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1554 , \oc8051_xiommu1/oc8051_page_table_i/n1555 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1556 , \oc8051_xiommu1/oc8051_page_table_i/n1557 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1558 , \oc8051_xiommu1/oc8051_page_table_i/n1559 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1560 , \oc8051_xiommu1/oc8051_page_table_i/n1561 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1562 , \oc8051_xiommu1/oc8051_page_table_i/n1563 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1564 , \oc8051_xiommu1/oc8051_page_table_i/n1565 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1566 , \oc8051_xiommu1/oc8051_page_table_i/n1567 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1568 , \oc8051_xiommu1/oc8051_page_table_i/n1569 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1570 , \oc8051_xiommu1/oc8051_page_table_i/n1571 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1572 , \oc8051_xiommu1/oc8051_page_table_i/n1573 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1574 , \oc8051_xiommu1/oc8051_page_table_i/n1575 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1576 , \oc8051_xiommu1/oc8051_page_table_i/n1577 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1578 , \oc8051_xiommu1/oc8051_page_table_i/n1579 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1580 , \oc8051_xiommu1/oc8051_page_table_i/n1581 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1582 , \oc8051_xiommu1/oc8051_page_table_i/n1583 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1584 , \oc8051_xiommu1/oc8051_page_table_i/n1585 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1586 , \oc8051_xiommu1/oc8051_page_table_i/n1587 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1588 , \oc8051_xiommu1/oc8051_page_table_i/n1589 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1590 , \oc8051_xiommu1/oc8051_page_table_i/n1591 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1592 , \oc8051_xiommu1/oc8051_page_table_i/n1593 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1594 , \oc8051_xiommu1/oc8051_page_table_i/n1595 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1596 , \oc8051_xiommu1/oc8051_page_table_i/n1597 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1598 , \oc8051_xiommu1/oc8051_page_table_i/n1599 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1600 , \oc8051_xiommu1/oc8051_page_table_i/n1601 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1602 , \oc8051_xiommu1/oc8051_page_table_i/n1603 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1604 , \oc8051_xiommu1/oc8051_page_table_i/n1605 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1606 , \oc8051_xiommu1/oc8051_page_table_i/n1607 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1608 , \oc8051_xiommu1/oc8051_page_table_i/n1609 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1610 , \oc8051_xiommu1/oc8051_page_table_i/n1611 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1612 , \oc8051_xiommu1/oc8051_page_table_i/n1613 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1614 , \oc8051_xiommu1/oc8051_page_table_i/n1615 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1616 , \oc8051_xiommu1/oc8051_page_table_i/n1617 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1618 , \oc8051_xiommu1/oc8051_page_table_i/n1619 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1620 , \oc8051_xiommu1/oc8051_page_table_i/n1621 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1622 , \oc8051_xiommu1/oc8051_page_table_i/n1623 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1624 , \oc8051_xiommu1/oc8051_page_table_i/n1625 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1626 , \oc8051_xiommu1/oc8051_page_table_i/n1627 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1628 , \oc8051_xiommu1/oc8051_page_table_i/n1629 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1630 , \oc8051_xiommu1/oc8051_page_table_i/n1631 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1632 , \oc8051_xiommu1/oc8051_page_table_i/n1633 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1634 , \oc8051_xiommu1/oc8051_page_table_i/n1635 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1636 , \oc8051_xiommu1/oc8051_page_table_i/n1637 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1638 , \oc8051_xiommu1/oc8051_page_table_i/n1639 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1640 , \oc8051_xiommu1/oc8051_page_table_i/n1641 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1642 , \oc8051_xiommu1/oc8051_page_table_i/n1643 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1644 , \oc8051_xiommu1/oc8051_page_table_i/n1645 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1646 , \oc8051_xiommu1/oc8051_page_table_i/n1647 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1648 , \oc8051_xiommu1/oc8051_page_table_i/n1649 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1650 , \oc8051_xiommu1/oc8051_page_table_i/n1651 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1652 , \oc8051_xiommu1/oc8051_page_table_i/n1653 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1654 , \oc8051_xiommu1/oc8051_page_table_i/n1655 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1656 , \oc8051_xiommu1/oc8051_page_table_i/n1657 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1658 , \oc8051_xiommu1/oc8051_page_table_i/n1659 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1660 , \oc8051_xiommu1/oc8051_page_table_i/n1661 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1662 , \oc8051_xiommu1/oc8051_page_table_i/n1663 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1664 , \oc8051_xiommu1/oc8051_page_table_i/n1665 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1666 , \oc8051_xiommu1/oc8051_page_table_i/n1667 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1668 , \oc8051_xiommu1/oc8051_page_table_i/n1669 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1670 , \oc8051_xiommu1/oc8051_page_table_i/n1671 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1672 , \oc8051_xiommu1/oc8051_page_table_i/n1673 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1674 , \oc8051_xiommu1/oc8051_page_table_i/n1675 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1676 , \oc8051_xiommu1/oc8051_page_table_i/n1677 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1678 , \oc8051_xiommu1/oc8051_page_table_i/n1679 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1680 , \oc8051_xiommu1/oc8051_page_table_i/n1681 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1682 , \oc8051_xiommu1/oc8051_page_table_i/n1683 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1684 , \oc8051_xiommu1/oc8051_page_table_i/n1685 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1686 , \oc8051_xiommu1/oc8051_page_table_i/n1687 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1688 , \oc8051_xiommu1/oc8051_page_table_i/n1689 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1690 , \oc8051_xiommu1/oc8051_page_table_i/n1691 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1692 , \oc8051_xiommu1/oc8051_page_table_i/n1693 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1694 , \oc8051_xiommu1/oc8051_page_table_i/n1695 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1696 , \oc8051_xiommu1/oc8051_page_table_i/n1697 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1698 , \oc8051_xiommu1/oc8051_page_table_i/n1699 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1700 , \oc8051_xiommu1/oc8051_page_table_i/n1701 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1702 , \oc8051_xiommu1/oc8051_page_table_i/n1703 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1704 , \oc8051_xiommu1/oc8051_page_table_i/n1705 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1706 , \oc8051_xiommu1/oc8051_page_table_i/n1707 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1708 , \oc8051_xiommu1/oc8051_page_table_i/n1709 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1710 , \oc8051_xiommu1/oc8051_page_table_i/n1711 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1712 , \oc8051_xiommu1/oc8051_page_table_i/n1713 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1714 , \oc8051_xiommu1/oc8051_page_table_i/n1715 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1716 , \oc8051_xiommu1/oc8051_page_table_i/n1717 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1718 , \oc8051_xiommu1/oc8051_page_table_i/n1719 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1720 , \oc8051_xiommu1/oc8051_page_table_i/n1721 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1722 , \oc8051_xiommu1/oc8051_page_table_i/n1723 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1724 , \oc8051_xiommu1/oc8051_page_table_i/n1725 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1726 , \oc8051_xiommu1/oc8051_page_table_i/n1727 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1728 , \oc8051_xiommu1/oc8051_page_table_i/n1729 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1730 , \oc8051_xiommu1/oc8051_page_table_i/n1731 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1732 , \oc8051_xiommu1/oc8051_page_table_i/n1733 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1734 , \oc8051_xiommu1/oc8051_page_table_i/n1735 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1736 , \oc8051_xiommu1/oc8051_page_table_i/n1737 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1738 , \oc8051_xiommu1/oc8051_page_table_i/n1739 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1740 , \oc8051_xiommu1/oc8051_page_table_i/n1741 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1742 , \oc8051_xiommu1/oc8051_page_table_i/n1743 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1744 , \oc8051_xiommu1/oc8051_page_table_i/n1745 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1746 , \oc8051_xiommu1/oc8051_page_table_i/n1747 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1748 , \oc8051_xiommu1/oc8051_page_table_i/n1749 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1750 , \oc8051_xiommu1/oc8051_page_table_i/n1751 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1752 , \oc8051_xiommu1/oc8051_page_table_i/n1753 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1754 , \oc8051_xiommu1/oc8051_page_table_i/n1755 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1756 , \oc8051_xiommu1/oc8051_page_table_i/n1757 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1758 , \oc8051_xiommu1/oc8051_page_table_i/n1759 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1760 , \oc8051_xiommu1/oc8051_page_table_i/n1761 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1762 , \oc8051_xiommu1/oc8051_page_table_i/n1763 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1764 , \oc8051_xiommu1/oc8051_page_table_i/n1765 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1766 , \oc8051_xiommu1/oc8051_page_table_i/n1767 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1768 , \oc8051_xiommu1/oc8051_page_table_i/n1769 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1770 , \oc8051_xiommu1/oc8051_page_table_i/n1771 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1772 , \oc8051_xiommu1/oc8051_page_table_i/n1773 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1774 , \oc8051_xiommu1/oc8051_page_table_i/n1775 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1776 , \oc8051_xiommu1/oc8051_page_table_i/n1777 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1778 , \oc8051_xiommu1/oc8051_page_table_i/n1779 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1780 , \oc8051_xiommu1/oc8051_page_table_i/n1781 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1782 , \oc8051_xiommu1/oc8051_page_table_i/n1783 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1784 , \oc8051_xiommu1/oc8051_page_table_i/n1785 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1786 , \oc8051_xiommu1/oc8051_page_table_i/n1787 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1788 , \oc8051_xiommu1/oc8051_page_table_i/n1789 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1790 , \oc8051_xiommu1/oc8051_page_table_i/n1791 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1792 , \oc8051_xiommu1/oc8051_page_table_i/n1793 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1794 , \oc8051_xiommu1/oc8051_page_table_i/n1795 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1796 , \oc8051_xiommu1/oc8051_page_table_i/n1797 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1798 , \oc8051_xiommu1/oc8051_page_table_i/n1799 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1800 , \oc8051_xiommu1/oc8051_page_table_i/n1801 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1802 , \oc8051_xiommu1/oc8051_page_table_i/n1803 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1804 , \oc8051_xiommu1/oc8051_page_table_i/n1805 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1806 , \oc8051_xiommu1/oc8051_page_table_i/n1807 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1808 , \oc8051_xiommu1/oc8051_page_table_i/n1809 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1810 , \oc8051_xiommu1/oc8051_page_table_i/n1811 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1812 , \oc8051_xiommu1/oc8051_page_table_i/n1813 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1814 , \oc8051_xiommu1/oc8051_page_table_i/n1815 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1816 , \oc8051_xiommu1/oc8051_page_table_i/n1817 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1818 , \oc8051_xiommu1/oc8051_page_table_i/n1819 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1820 , \oc8051_xiommu1/oc8051_page_table_i/n1821 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1822 , \oc8051_xiommu1/oc8051_page_table_i/n1823 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1824 , \oc8051_xiommu1/oc8051_page_table_i/n1825 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1826 , \oc8051_xiommu1/oc8051_page_table_i/n1827 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1828 , \oc8051_xiommu1/oc8051_page_table_i/n1829 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1830 , \oc8051_xiommu1/oc8051_page_table_i/n1831 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1832 , \oc8051_xiommu1/oc8051_page_table_i/n1833 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1834 , \oc8051_xiommu1/oc8051_page_table_i/n1835 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1836 , \oc8051_xiommu1/oc8051_page_table_i/n1837 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1838 , \oc8051_xiommu1/oc8051_page_table_i/n1839 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1840 , \oc8051_xiommu1/oc8051_page_table_i/n1841 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1842 , \oc8051_xiommu1/oc8051_page_table_i/n1843 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1844 , \oc8051_xiommu1/oc8051_page_table_i/n1845 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1846 , \oc8051_xiommu1/oc8051_page_table_i/n1847 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1848 , \oc8051_xiommu1/oc8051_page_table_i/n1849 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1850 , \oc8051_xiommu1/oc8051_page_table_i/n1851 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1852 , \oc8051_xiommu1/oc8051_page_table_i/n1853 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1854 , \oc8051_xiommu1/oc8051_page_table_i/n1855 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1856 , \oc8051_xiommu1/oc8051_page_table_i/n1857 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1858 , \oc8051_xiommu1/oc8051_page_table_i/n1859 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1860 , \oc8051_xiommu1/oc8051_page_table_i/n1861 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1862 , \oc8051_xiommu1/oc8051_page_table_i/n1863 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1864 , \oc8051_xiommu1/oc8051_page_table_i/n1865 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1866 , \oc8051_xiommu1/oc8051_page_table_i/n1867 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1868 , \oc8051_xiommu1/oc8051_page_table_i/n1869 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1870 , \oc8051_xiommu1/oc8051_page_table_i/n1871 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1872 , \oc8051_xiommu1/oc8051_page_table_i/n1873 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1874 , \oc8051_xiommu1/oc8051_page_table_i/n1875 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1876 , \oc8051_xiommu1/oc8051_page_table_i/n1877 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1878 , \oc8051_xiommu1/oc8051_page_table_i/n1879 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1880 , \oc8051_xiommu1/oc8051_page_table_i/n1881 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1882 , \oc8051_xiommu1/oc8051_page_table_i/n1883 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1884 , \oc8051_xiommu1/oc8051_page_table_i/n1885 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1886 , \oc8051_xiommu1/oc8051_page_table_i/n1887 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1888 , \oc8051_xiommu1/oc8051_page_table_i/n1889 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1890 , \oc8051_xiommu1/oc8051_page_table_i/n1891 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1892 , \oc8051_xiommu1/oc8051_page_table_i/n1893 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1894 , \oc8051_xiommu1/oc8051_page_table_i/n1895 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1896 , \oc8051_xiommu1/oc8051_page_table_i/n1897 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1898 , \oc8051_xiommu1/oc8051_page_table_i/n1899 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1900 , \oc8051_xiommu1/oc8051_page_table_i/n1901 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1902 , \oc8051_xiommu1/oc8051_page_table_i/n1903 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1904 , \oc8051_xiommu1/oc8051_page_table_i/n1905 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1906 , \oc8051_xiommu1/oc8051_page_table_i/n1907 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1908 , \oc8051_xiommu1/oc8051_page_table_i/n1909 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1910 , \oc8051_xiommu1/oc8051_page_table_i/n1911 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1912 , \oc8051_xiommu1/oc8051_page_table_i/n1913 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1914 , \oc8051_xiommu1/oc8051_page_table_i/n1915 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1916 , \oc8051_xiommu1/oc8051_page_table_i/n1917 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1918 , \oc8051_xiommu1/oc8051_page_table_i/n1919 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1920 , \oc8051_xiommu1/oc8051_page_table_i/n1921 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1922 , \oc8051_xiommu1/oc8051_page_table_i/n1923 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1924 , \oc8051_xiommu1/oc8051_page_table_i/n1925 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1926 , \oc8051_xiommu1/oc8051_page_table_i/n1927 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1928 , \oc8051_xiommu1/oc8051_page_table_i/n1929 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1930 , \oc8051_xiommu1/oc8051_page_table_i/n1931 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1932 , \oc8051_xiommu1/oc8051_page_table_i/n1933 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1934 , \oc8051_xiommu1/oc8051_page_table_i/n1935 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1936 , \oc8051_xiommu1/oc8051_page_table_i/n1937 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1938 , \oc8051_xiommu1/oc8051_page_table_i/n1939 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1940 , \oc8051_xiommu1/oc8051_page_table_i/n1941 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1942 , \oc8051_xiommu1/oc8051_page_table_i/n1943 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1944 , \oc8051_xiommu1/oc8051_page_table_i/n1945 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1946 , \oc8051_xiommu1/oc8051_page_table_i/n1947 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1948 , \oc8051_xiommu1/oc8051_page_table_i/n1949 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1950 , \oc8051_xiommu1/oc8051_page_table_i/n1951 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1952 , \oc8051_xiommu1/oc8051_page_table_i/n1953 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1954 , \oc8051_xiommu1/oc8051_page_table_i/n1955 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1956 , \oc8051_xiommu1/oc8051_page_table_i/n1957 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1958 , \oc8051_xiommu1/oc8051_page_table_i/n1959 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1960 , \oc8051_xiommu1/oc8051_page_table_i/n1961 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1962 , \oc8051_xiommu1/oc8051_page_table_i/n1963 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1964 , \oc8051_xiommu1/oc8051_page_table_i/n1965 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1966 , \oc8051_xiommu1/oc8051_page_table_i/n1967 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1968 , \oc8051_xiommu1/oc8051_page_table_i/n1969 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1970 , \oc8051_xiommu1/oc8051_page_table_i/n1971 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1972 , \oc8051_xiommu1/oc8051_page_table_i/n1973 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1974 , \oc8051_xiommu1/oc8051_page_table_i/n1975 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1976 , \oc8051_xiommu1/oc8051_page_table_i/n1977 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1978 , \oc8051_xiommu1/oc8051_page_table_i/n1979 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1980 , \oc8051_xiommu1/oc8051_page_table_i/n1981 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1982 , \oc8051_xiommu1/oc8051_page_table_i/n1983 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1984 , \oc8051_xiommu1/oc8051_page_table_i/n1985 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1986 , \oc8051_xiommu1/oc8051_page_table_i/n1987 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1988 , \oc8051_xiommu1/oc8051_page_table_i/n1989 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1990 , \oc8051_xiommu1/oc8051_page_table_i/n1991 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1992 , \oc8051_xiommu1/oc8051_page_table_i/n1993 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1994 , \oc8051_xiommu1/oc8051_page_table_i/n1995 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1996 , \oc8051_xiommu1/oc8051_page_table_i/n1997 , 
        \oc8051_xiommu1/oc8051_page_table_i/n1998 , \oc8051_xiommu1/oc8051_page_table_i/n1999 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2000 , \oc8051_xiommu1/oc8051_page_table_i/n2001 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2002 , \oc8051_xiommu1/oc8051_page_table_i/n2003 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2004 , \oc8051_xiommu1/oc8051_page_table_i/n2005 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2006 , \oc8051_xiommu1/oc8051_page_table_i/n2007 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2008 , \oc8051_xiommu1/oc8051_page_table_i/n2009 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2010 , \oc8051_xiommu1/oc8051_page_table_i/n2011 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2012 , \oc8051_xiommu1/oc8051_page_table_i/n2013 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2014 , \oc8051_xiommu1/oc8051_page_table_i/n2015 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2016 , \oc8051_xiommu1/oc8051_page_table_i/n2017 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2018 , \oc8051_xiommu1/oc8051_page_table_i/n2531 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2532 , \oc8051_xiommu1/oc8051_page_table_i/n2534 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2535 , \oc8051_xiommu1/oc8051_page_table_i/n2536 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2542 , \oc8051_xiommu1/oc8051_page_table_i/n2567 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2568 , \oc8051_xiommu1/oc8051_page_table_i/n2569 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2570 , \oc8051_xiommu1/oc8051_page_table_i/n2571 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2572 , \oc8051_xiommu1/oc8051_page_table_i/n2573 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2574 , \oc8051_xiommu1/oc8051_page_table_i/n2575 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2576 , \oc8051_xiommu1/oc8051_page_table_i/n2577 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2578 , \oc8051_xiommu1/oc8051_page_table_i/n2579 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2580 , \oc8051_xiommu1/oc8051_page_table_i/n2581 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2582 , \oc8051_xiommu1/oc8051_page_table_i/n2583 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2584 , \oc8051_xiommu1/oc8051_page_table_i/n2585 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2586 , \oc8051_xiommu1/oc8051_page_table_i/n2587 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2588 , \oc8051_xiommu1/oc8051_page_table_i/n2589 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2590 , \oc8051_xiommu1/oc8051_page_table_i/n2591 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2592 , \oc8051_xiommu1/oc8051_page_table_i/n2593 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2594 , \oc8051_xiommu1/oc8051_page_table_i/n2595 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2596 , \oc8051_xiommu1/oc8051_page_table_i/n2597 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2598 , \oc8051_xiommu1/oc8051_page_table_i/n2610 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2612 , \oc8051_xiommu1/oc8051_page_table_i/n2613 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2614 , \oc8051_xiommu1/oc8051_page_table_i/n2615 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2616 , \oc8051_xiommu1/oc8051_page_table_i/n2617 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2618 , \oc8051_xiommu1/oc8051_page_table_i/n2619 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2620 , \oc8051_xiommu1/oc8051_page_table_i/n2621 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2622 , \oc8051_xiommu1/oc8051_page_table_i/n2623 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2624 , \oc8051_xiommu1/oc8051_page_table_i/n2625 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2626 , \oc8051_xiommu1/oc8051_page_table_i/n2627 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2628 , \oc8051_xiommu1/oc8051_page_table_i/n2629 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2630 , \oc8051_xiommu1/oc8051_page_table_i/n2631 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2632 , \oc8051_xiommu1/oc8051_page_table_i/n2633 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2634 , \oc8051_xiommu1/oc8051_page_table_i/n2635 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2636 , \oc8051_xiommu1/oc8051_page_table_i/n2637 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2638 , \oc8051_xiommu1/oc8051_page_table_i/n2639 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2640 , \oc8051_xiommu1/oc8051_page_table_i/n2641 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2642 , \oc8051_xiommu1/oc8051_page_table_i/n2643 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2644 , \oc8051_xiommu1/oc8051_page_table_i/n2645 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2646 , \oc8051_xiommu1/oc8051_page_table_i/n2647 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2648 , \oc8051_xiommu1/oc8051_page_table_i/n2649 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2650 , \oc8051_xiommu1/oc8051_page_table_i/n2651 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2652 , \oc8051_xiommu1/oc8051_page_table_i/n2653 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2654 , \oc8051_xiommu1/oc8051_page_table_i/n2655 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2656 , \oc8051_xiommu1/oc8051_page_table_i/n2657 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2658 , \oc8051_xiommu1/oc8051_page_table_i/n2659 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2660 , \oc8051_xiommu1/oc8051_page_table_i/n2661 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2662 , \oc8051_xiommu1/oc8051_page_table_i/n2663 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2664 , \oc8051_xiommu1/oc8051_page_table_i/n2665 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2666 , \oc8051_xiommu1/oc8051_page_table_i/n2667 , 
        \oc8051_xiommu1/oc8051_page_table_i/n2668 , \oc8051_xiommu1/aes_top_i/LessThan_3/n2 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n4 , \oc8051_xiommu1/aes_top_i/LessThan_3/n6 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n8 , \oc8051_xiommu1/aes_top_i/LessThan_3/n10 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n12 , \oc8051_xiommu1/aes_top_i/LessThan_3/n14 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n16 , \oc8051_xiommu1/aes_top_i/LessThan_3/n18 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n20 , \oc8051_xiommu1/aes_top_i/LessThan_3/n22 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n24 , \oc8051_xiommu1/aes_top_i/LessThan_3/n26 , 
        \oc8051_xiommu1/aes_top_i/LessThan_3/n28 , \oc8051_xiommu1/aes_top_i/LessThan_3/n30 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n2 , \oc8051_xiommu1/aes_top_i/LessThan_4/n4 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n6 , \oc8051_xiommu1/aes_top_i/LessThan_4/n8 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n10 , \oc8051_xiommu1/aes_top_i/LessThan_4/n12 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n14 , \oc8051_xiommu1/aes_top_i/LessThan_4/n16 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n18 , \oc8051_xiommu1/aes_top_i/LessThan_4/n20 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n22 , \oc8051_xiommu1/aes_top_i/LessThan_4/n24 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n26 , \oc8051_xiommu1/aes_top_i/LessThan_4/n28 , 
        \oc8051_xiommu1/aes_top_i/LessThan_4/n30 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n4 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n8 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n9 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n12 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n13 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n15 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n12 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n14 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n15 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n4 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n8 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n9 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n12 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n13 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n15 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n12 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n14 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n12 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n14 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n4 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n8 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n9 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_144/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_146/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_148/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_151/n1 , \oc8051_xiommu1/aes_top_i/add_163/n2 , 
        \oc8051_xiommu1/aes_top_i/add_163/n4 , \oc8051_xiommu1/aes_top_i/add_163/n6 , 
        \oc8051_xiommu1/aes_top_i/add_163/n8 , \oc8051_xiommu1/aes_top_i/add_163/n10 , 
        \oc8051_xiommu1/aes_top_i/add_163/n12 , \oc8051_xiommu1/aes_top_i/add_163/n14 , 
        \oc8051_xiommu1/aes_top_i/add_163/n16 , \oc8051_xiommu1/aes_top_i/add_163/n18 , 
        \oc8051_xiommu1/aes_top_i/add_163/n20 , \oc8051_xiommu1/aes_top_i/add_163/n22 , 
        \oc8051_xiommu1/aes_top_i/add_163/cout , \oc8051_xiommu1/aes_top_i/add_194/n2 , 
        \oc8051_xiommu1/aes_top_i/add_194/n4 , \oc8051_xiommu1/aes_top_i/add_194/n6 , 
        \oc8051_xiommu1/aes_top_i/add_194/n8 , \oc8051_xiommu1/aes_top_i/add_194/n10 , 
        \oc8051_xiommu1/aes_top_i/add_194/n12 , \oc8051_xiommu1/aes_top_i/add_194/n14 , 
        \oc8051_xiommu1/aes_top_i/add_194/n16 , \oc8051_xiommu1/aes_top_i/add_194/n18 , 
        \oc8051_xiommu1/aes_top_i/add_194/n20 , \oc8051_xiommu1/aes_top_i/add_194/n22 , 
        \oc8051_xiommu1/aes_top_i/add_194/cout , \oc8051_xiommu1/aes_top_i/add_225/n2 , 
        \oc8051_xiommu1/aes_top_i/add_225/n4 , \oc8051_xiommu1/aes_top_i/add_225/n6 , 
        \oc8051_xiommu1/aes_top_i/add_225/cout , \oc8051_xiommu1/aes_top_i/reduce_nor_240/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_240/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_240/n3 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n2 , \oc8051_xiommu1/aes_top_i/LessThan_243/n4 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n6 , \oc8051_xiommu1/aes_top_i/LessThan_243/n8 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n10 , \oc8051_xiommu1/aes_top_i/LessThan_243/n12 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n14 , \oc8051_xiommu1/aes_top_i/LessThan_243/n16 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n18 , \oc8051_xiommu1/aes_top_i/LessThan_243/n20 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n22 , \oc8051_xiommu1/aes_top_i/LessThan_243/n24 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n26 , \oc8051_xiommu1/aes_top_i/LessThan_243/n28 , 
        \oc8051_xiommu1/aes_top_i/LessThan_243/n30 , \oc8051_xiommu1/aes_top_i/add_245/n2 , 
        \oc8051_xiommu1/aes_top_i/add_245/n4 , \oc8051_xiommu1/aes_top_i/add_245/n6 , 
        \oc8051_xiommu1/aes_top_i/add_245/n8 , \oc8051_xiommu1/aes_top_i/add_245/n10 , 
        \oc8051_xiommu1/aes_top_i/add_245/n12 , \oc8051_xiommu1/aes_top_i/add_245/n14 , 
        \oc8051_xiommu1/aes_top_i/add_245/n16 , \oc8051_xiommu1/aes_top_i/add_245/n18 , 
        \oc8051_xiommu1/aes_top_i/add_245/n20 , \oc8051_xiommu1/aes_top_i/add_245/n22 , 
        \oc8051_xiommu1/aes_top_i/add_245/n24 , \oc8051_xiommu1/aes_top_i/add_245/n26 , 
        \oc8051_xiommu1/aes_top_i/add_245/n28 , \oc8051_xiommu1/aes_top_i/add_245/n30 , 
        \oc8051_xiommu1/aes_top_i/add_245/cout , \oc8051_xiommu1/aes_top_i/add_246/n2 , 
        \oc8051_xiommu1/aes_top_i/add_246/n4 , \oc8051_xiommu1/aes_top_i/add_246/n6 , 
        \oc8051_xiommu1/aes_top_i/add_246/n8 , \oc8051_xiommu1/aes_top_i/add_246/n10 , 
        \oc8051_xiommu1/aes_top_i/add_246/n12 , \oc8051_xiommu1/aes_top_i/add_246/n14 , 
        \oc8051_xiommu1/aes_top_i/add_246/n16 , \oc8051_xiommu1/aes_top_i/add_246/n18 , 
        \oc8051_xiommu1/aes_top_i/add_246/n20 , \oc8051_xiommu1/aes_top_i/add_246/n22 , 
        \oc8051_xiommu1/aes_top_i/add_246/n24 , \oc8051_xiommu1/aes_top_i/add_246/n26 , 
        \oc8051_xiommu1/aes_top_i/add_246/n28 , \oc8051_xiommu1/aes_top_i/add_246/n30 , 
        \oc8051_xiommu1/aes_top_i/add_246/cout , \oc8051_xiommu1/aes_top_i/reduce_nor_265/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_265/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_265/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_276/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_276/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_276/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_287/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_287/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_287/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_299/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_299/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_299/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_310/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_310/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_310/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_322/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_322/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_322/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_334/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_334/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_334/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_347/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_347/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_347/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_358/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_358/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_358/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_370/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_370/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_370/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_382/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_382/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_382/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_395/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_395/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_395/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_407/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_407/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_407/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_420/n1 , \oc8051_xiommu1/aes_top_i/reduce_nor_420/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_420/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_433/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_433/n2 , \oc8051_xiommu1/aes_top_i/reduce_nor_433/n3 , 
        \oc8051_xiommu1/aes_top_i/add_457/n2 , \oc8051_xiommu1/aes_top_i/add_457/n4 , 
        \oc8051_xiommu1/aes_top_i/add_457/n6 , \oc8051_xiommu1/aes_top_i/add_457/n8 , 
        \oc8051_xiommu1/aes_top_i/add_457/n10 , \oc8051_xiommu1/aes_top_i/add_457/n12 , 
        \oc8051_xiommu1/aes_top_i/add_457/n14 , \oc8051_xiommu1/aes_top_i/add_457/n16 , 
        \oc8051_xiommu1/aes_top_i/add_457/n18 , \oc8051_xiommu1/aes_top_i/add_457/n20 , 
        \oc8051_xiommu1/aes_top_i/add_457/n22 , \oc8051_xiommu1/aes_top_i/add_457/n24 , 
        \oc8051_xiommu1/aes_top_i/add_457/n26 , \oc8051_xiommu1/aes_top_i/add_457/n28 , 
        \oc8051_xiommu1/aes_top_i/add_457/n30 , \oc8051_xiommu1/aes_top_i/add_457/n32 , 
        \oc8051_xiommu1/aes_top_i/add_457/n34 , \oc8051_xiommu1/aes_top_i/add_457/n36 , 
        \oc8051_xiommu1/aes_top_i/add_457/n38 , \oc8051_xiommu1/aes_top_i/add_457/n40 , 
        \oc8051_xiommu1/aes_top_i/add_457/n42 , \oc8051_xiommu1/aes_top_i/add_457/n44 , 
        \oc8051_xiommu1/aes_top_i/add_457/n46 , \oc8051_xiommu1/aes_top_i/add_457/n48 , 
        \oc8051_xiommu1/aes_top_i/add_457/n50 , \oc8051_xiommu1/aes_top_i/add_457/n52 , 
        \oc8051_xiommu1/aes_top_i/add_457/n54 , \oc8051_xiommu1/aes_top_i/add_457/n56 , 
        \oc8051_xiommu1/aes_top_i/add_457/n58 , \oc8051_xiommu1/aes_top_i/add_457/n60 , 
        \oc8051_xiommu1/aes_top_i/add_457/n62 , \oc8051_xiommu1/aes_top_i/add_457/n64 , 
        \oc8051_xiommu1/aes_top_i/add_457/n66 , \oc8051_xiommu1/aes_top_i/add_457/n68 , 
        \oc8051_xiommu1/aes_top_i/add_457/n70 , \oc8051_xiommu1/aes_top_i/add_457/n72 , 
        \oc8051_xiommu1/aes_top_i/add_457/n74 , \oc8051_xiommu1/aes_top_i/add_457/n76 , 
        \oc8051_xiommu1/aes_top_i/add_457/n78 , \oc8051_xiommu1/aes_top_i/add_457/n80 , 
        \oc8051_xiommu1/aes_top_i/add_457/n82 , \oc8051_xiommu1/aes_top_i/add_457/n84 , 
        \oc8051_xiommu1/aes_top_i/add_457/n86 , \oc8051_xiommu1/aes_top_i/add_457/n88 , 
        \oc8051_xiommu1/aes_top_i/add_457/n90 , \oc8051_xiommu1/aes_top_i/add_457/n92 , 
        \oc8051_xiommu1/aes_top_i/add_457/n94 , \oc8051_xiommu1/aes_top_i/add_457/n96 , 
        \oc8051_xiommu1/aes_top_i/add_457/n98 , \oc8051_xiommu1/aes_top_i/add_457/n100 , 
        \oc8051_xiommu1/aes_top_i/add_457/n102 , \oc8051_xiommu1/aes_top_i/add_457/n104 , 
        \oc8051_xiommu1/aes_top_i/add_457/n106 , \oc8051_xiommu1/aes_top_i/add_457/n108 , 
        \oc8051_xiommu1/aes_top_i/add_457/n110 , \oc8051_xiommu1/aes_top_i/add_457/n112 , 
        \oc8051_xiommu1/aes_top_i/add_457/n114 , \oc8051_xiommu1/aes_top_i/add_457/n116 , 
        \oc8051_xiommu1/aes_top_i/add_457/n118 , \oc8051_xiommu1/aes_top_i/add_457/n120 , 
        \oc8051_xiommu1/aes_top_i/add_457/n122 , \oc8051_xiommu1/aes_top_i/add_457/n124 , 
        \oc8051_xiommu1/aes_top_i/add_457/n126 , \oc8051_xiommu1/aes_top_i/add_457/n128 , 
        \oc8051_xiommu1/aes_top_i/add_457/n130 , \oc8051_xiommu1/aes_top_i/add_457/n132 , 
        \oc8051_xiommu1/aes_top_i/add_457/n134 , \oc8051_xiommu1/aes_top_i/add_457/n136 , 
        \oc8051_xiommu1/aes_top_i/add_457/n138 , \oc8051_xiommu1/aes_top_i/add_457/n140 , 
        \oc8051_xiommu1/aes_top_i/add_457/n142 , \oc8051_xiommu1/aes_top_i/add_457/n144 , 
        \oc8051_xiommu1/aes_top_i/add_457/n146 , \oc8051_xiommu1/aes_top_i/add_457/n148 , 
        \oc8051_xiommu1/aes_top_i/add_457/n150 , \oc8051_xiommu1/aes_top_i/add_457/n152 , 
        \oc8051_xiommu1/aes_top_i/add_457/n154 , \oc8051_xiommu1/aes_top_i/add_457/n156 , 
        \oc8051_xiommu1/aes_top_i/add_457/n158 , \oc8051_xiommu1/aes_top_i/add_457/n160 , 
        \oc8051_xiommu1/aes_top_i/add_457/n162 , \oc8051_xiommu1/aes_top_i/add_457/n164 , 
        \oc8051_xiommu1/aes_top_i/add_457/n166 , \oc8051_xiommu1/aes_top_i/add_457/n168 , 
        \oc8051_xiommu1/aes_top_i/add_457/n170 , \oc8051_xiommu1/aes_top_i/add_457/n172 , 
        \oc8051_xiommu1/aes_top_i/add_457/n174 , \oc8051_xiommu1/aes_top_i/add_457/n176 , 
        \oc8051_xiommu1/aes_top_i/add_457/n178 , \oc8051_xiommu1/aes_top_i/add_457/n180 , 
        \oc8051_xiommu1/aes_top_i/add_457/n182 , \oc8051_xiommu1/aes_top_i/add_457/n184 , 
        \oc8051_xiommu1/aes_top_i/add_457/n186 , \oc8051_xiommu1/aes_top_i/add_457/n188 , 
        \oc8051_xiommu1/aes_top_i/add_457/n190 , \oc8051_xiommu1/aes_top_i/add_457/n192 , 
        \oc8051_xiommu1/aes_top_i/add_457/n194 , \oc8051_xiommu1/aes_top_i/add_457/n196 , 
        \oc8051_xiommu1/aes_top_i/add_457/n198 , \oc8051_xiommu1/aes_top_i/add_457/n200 , 
        \oc8051_xiommu1/aes_top_i/add_457/n202 , \oc8051_xiommu1/aes_top_i/add_457/n204 , 
        \oc8051_xiommu1/aes_top_i/add_457/n206 , \oc8051_xiommu1/aes_top_i/add_457/n208 , 
        \oc8051_xiommu1/aes_top_i/add_457/n210 , \oc8051_xiommu1/aes_top_i/add_457/n212 , 
        \oc8051_xiommu1/aes_top_i/add_457/n214 , \oc8051_xiommu1/aes_top_i/add_457/n216 , 
        \oc8051_xiommu1/aes_top_i/add_457/n218 , \oc8051_xiommu1/aes_top_i/add_457/n220 , 
        \oc8051_xiommu1/aes_top_i/add_457/n222 , \oc8051_xiommu1/aes_top_i/add_457/n224 , 
        \oc8051_xiommu1/aes_top_i/add_457/n226 , \oc8051_xiommu1/aes_top_i/add_457/n228 , 
        \oc8051_xiommu1/aes_top_i/add_457/n230 , \oc8051_xiommu1/aes_top_i/add_457/n232 , 
        \oc8051_xiommu1/aes_top_i/add_457/n234 , \oc8051_xiommu1/aes_top_i/add_457/n236 , 
        \oc8051_xiommu1/aes_top_i/add_457/n238 , \oc8051_xiommu1/aes_top_i/add_457/n240 , 
        \oc8051_xiommu1/aes_top_i/add_457/n242 , \oc8051_xiommu1/aes_top_i/add_457/n244 , 
        \oc8051_xiommu1/aes_top_i/add_457/n246 , \oc8051_xiommu1/aes_top_i/add_457/n248 , 
        \oc8051_xiommu1/aes_top_i/add_457/n250 , \oc8051_xiommu1/aes_top_i/add_457/n252 , 
        \oc8051_xiommu1/aes_top_i/add_457/n254 , \oc8051_xiommu1/aes_top_i/add_457/cout , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n2 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n2 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n2 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n2 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n2 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n6 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n10 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n14 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n18 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n22 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n26 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n30 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n4 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n8 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n12 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n16 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n20 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n24 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n28 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n2 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n6 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n10 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n14 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n18 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n22 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n26 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n30 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n4 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n8 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n12 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n16 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n20 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n24 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n28 , \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n1 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n5 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n9 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n11 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n2 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n4 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n5 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n8 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n9 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n12 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n1 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n5 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n9 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n11 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n2 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n4 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n5 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n8 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n9 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n12 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n1 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n5 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n9 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n11 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n2 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n4 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n5 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n8 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n9 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n12 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n1 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n2 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n3 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n5 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n7 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n9 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n11 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n13 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n15 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n17 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n19 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n21 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n23 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n25 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n27 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n29 , \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n3 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n8 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n9 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n10 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n12 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n14 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n16 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n18 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n20 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n21 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n22 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n23 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n24 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n25 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n26 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n27 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n28 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n29 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n30 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n31 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n32 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n33 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n34 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n35 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n36 , \oc8051_xiommu1/oc8051_page_table_i/reduce_or_2475/n1 ;
    
    assign _cvpt_914 = rst;   // oc8051_tb.v(112)
    assign _cvpt_1 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_2 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_3 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_4 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_5 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_6 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_7 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_8 = _cvpt_0;   // oc8051_tb.v(104)
    assign _cvpt_10 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_12 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_13 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_14 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_15 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_16 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_17 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_18 = _cvpt_11;   // oc8051_tb.v(104)
    assign _cvpt_20 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_21 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_22 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_23 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_24 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_25 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_26 = _cvpt_19;   // oc8051_tb.v(104)
    assign _cvpt_27 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_28 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_29 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_30 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_31 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_32 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_33 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_34 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_35 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_36 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_37 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_38 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_39 = _cvpt_9;   // oc8051_tb.v(104)
    assign _cvpt_42 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_43 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_44 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_45 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_46 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_47 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_48 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_49 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_50 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_51 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_52 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_53 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_54 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_55 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_56 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_57 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_58 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_59 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_60 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_61 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_62 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_63 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_64 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_65 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_66 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_67 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_68 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_69 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_70 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_71 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_72 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_73 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_74 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_76 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_77 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_78 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_79 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_80 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_81 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_82 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_83 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_84 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_85 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_86 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_87 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_88 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_89 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_90 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_91 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_92 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_93 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_94 = _cvpt_75;   // oc8051_tb.v(104)
    assign _cvpt_96 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_97 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_98 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_99 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_100 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_101 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_102 = _cvpt_95;   // oc8051_tb.v(104)
    assign _cvpt_105 = _cvpt_104;   // oc8051_tb.v(104)
    assign _cvpt_107 = _cvpt_106;   // oc8051_tb.v(104)
    assign _cvpt_109 = _cvpt_108;   // oc8051_tb.v(104)
    assign _cvpt_110 = _cvpt_108;   // oc8051_tb.v(104)
    assign _cvpt_112 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_113 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_114 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_115 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_116 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_117 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_118 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_120 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_121 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_122 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_123 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_124 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_125 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_126 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_128 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_129 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_130 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_131 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_132 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_133 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_134 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_136 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_137 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_138 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_139 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_140 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_141 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_142 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_144 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_145 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_146 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_147 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_148 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_149 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_150 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_152 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_153 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_154 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_155 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_156 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_157 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_158 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_159 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_160 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_161 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_162 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_163 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_164 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_165 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_166 = _cvpt_111;   // oc8051_tb.v(104)
    assign _cvpt_167 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_168 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_169 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_170 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_171 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_172 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_173 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_174 = _cvpt_119;   // oc8051_tb.v(104)
    assign _cvpt_175 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_176 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_177 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_178 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_179 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_180 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_181 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_182 = _cvpt_127;   // oc8051_tb.v(104)
    assign _cvpt_183 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_184 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_185 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_186 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_187 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_188 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_189 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_190 = _cvpt_135;   // oc8051_tb.v(104)
    assign _cvpt_191 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_192 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_193 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_194 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_195 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_196 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_197 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_198 = _cvpt_143;   // oc8051_tb.v(104)
    assign _cvpt_199 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_200 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_201 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_202 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_203 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_204 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_205 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_206 = _cvpt_151;   // oc8051_tb.v(104)
    assign _cvpt_207 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_209 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_210 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_211 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_212 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_213 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_214 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_215 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_216 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_217 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_218 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_219 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_220 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_221 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_222 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_223 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_224 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_225 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_226 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_227 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_228 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_229 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_230 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_231 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_232 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_233 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_234 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_235 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_236 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_237 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_238 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_239 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_240 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_241 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_242 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_243 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_244 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_245 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_246 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_247 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_248 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_249 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_250 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_251 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_252 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_253 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_254 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_255 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_256 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_257 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_258 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_259 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_260 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_261 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_262 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_263 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_264 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_265 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_266 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_267 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_268 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_269 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_270 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_271 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_272 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_273 = _cvpt_40;   // oc8051_tb.v(104)
    assign _cvpt_274 = _cvpt_208;   // oc8051_tb.v(104)
    assign _cvpt_275 = _cvpt_104;   // oc8051_tb.v(104)
    assign _cvpt_277 = _cvpt_104;   // oc8051_tb.v(104)
    assign _cvpt_278 = _cvpt_276;   // oc8051_tb.v(104)
    assign _cvpt_280 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_281 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_282 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_283 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_284 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_285 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_286 = _cvpt_279;   // oc8051_tb.v(104)
    assign _cvpt_288 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_289 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_290 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_291 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_292 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_293 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_294 = _cvpt_287;   // oc8051_tb.v(104)
    assign _cvpt_296 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_297 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_298 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_299 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_300 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_301 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_302 = _cvpt_295;   // oc8051_tb.v(104)
    assign _cvpt_304 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_305 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_306 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_307 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_308 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_309 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_310 = _cvpt_303;   // oc8051_tb.v(104)
    assign _cvpt_312 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_313 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_314 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_315 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_316 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_317 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_318 = _cvpt_311;   // oc8051_tb.v(104)
    assign _cvpt_320 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_321 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_322 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_323 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_324 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_325 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_326 = _cvpt_319;   // oc8051_tb.v(104)
    assign _cvpt_328 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_329 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_330 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_331 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_332 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_333 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_334 = _cvpt_327;   // oc8051_tb.v(104)
    assign _cvpt_337 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_338 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_339 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_340 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_341 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_342 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_343 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_344 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_345 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_346 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_347 = _cvpt_336;   // oc8051_tb.v(104)
    assign _cvpt_349 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_350 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_351 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_352 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_353 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_354 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_355 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_356 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_357 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_358 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_359 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_360 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_361 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_362 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_363 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_365 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_366 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_367 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_368 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_369 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_370 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_371 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_372 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_373 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_374 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_375 = _cvpt_364;   // oc8051_tb.v(104)
    assign _cvpt_376 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_377 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_378 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_379 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_380 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_381 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_382 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_383 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_384 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_385 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_386 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_387 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_388 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_389 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_390 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_391 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_393 = _cvpt_392;   // oc8051_tb.v(104)
    assign _cvpt_394 = _cvpt_392;   // oc8051_tb.v(104)
    assign _cvpt_395 = _cvpt_392;   // oc8051_tb.v(104)
    assign _cvpt_396 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_397 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_398 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_399 = _cvpt_348;   // oc8051_tb.v(104)
    assign _cvpt_401 = _cvpt_400;   // oc8051_tb.v(104)
    assign _cvpt_403 = _cvpt_402;   // oc8051_tb.v(104)
    assign _cvpt_405 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_407 = _cvpt_406;   // oc8051_tb.v(104)
    assign _cvpt_409 = _cvpt_408;   // oc8051_tb.v(104)
    assign _cvpt_411 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_412 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_413 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_414 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_415 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_416 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_417 = _cvpt_410;   // oc8051_tb.v(104)
    assign _cvpt_419 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_420 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_421 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_422 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_423 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_424 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_425 = _cvpt_418;   // oc8051_tb.v(104)
    assign _cvpt_427 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_428 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_429 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_430 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_431 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_432 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_433 = _cvpt_426;   // oc8051_tb.v(104)
    assign _cvpt_435 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_436 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_437 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_438 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_439 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_440 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_441 = _cvpt_434;   // oc8051_tb.v(104)
    assign _cvpt_443 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_444 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_445 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_446 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_447 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_448 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_449 = _cvpt_442;   // oc8051_tb.v(104)
    assign _cvpt_451 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_452 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_453 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_454 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_455 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_456 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_457 = _cvpt_450;   // oc8051_tb.v(104)
    assign _cvpt_459 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_460 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_461 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_462 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_463 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_464 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_465 = _cvpt_458;   // oc8051_tb.v(104)
    assign _cvpt_467 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_468 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_469 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_470 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_471 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_472 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_473 = _cvpt_466;   // oc8051_tb.v(104)
    assign _cvpt_475 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_476 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_477 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_478 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_479 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_480 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_481 = _cvpt_474;   // oc8051_tb.v(104)
    assign _cvpt_483 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_484 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_485 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_486 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_487 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_488 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_489 = _cvpt_482;   // oc8051_tb.v(104)
    assign _cvpt_491 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_492 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_493 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_494 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_495 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_496 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_497 = _cvpt_490;   // oc8051_tb.v(104)
    assign _cvpt_499 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_500 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_501 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_502 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_503 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_504 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_505 = _cvpt_498;   // oc8051_tb.v(104)
    assign _cvpt_507 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_508 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_509 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_510 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_511 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_512 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_513 = _cvpt_506;   // oc8051_tb.v(104)
    assign _cvpt_515 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_516 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_517 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_518 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_519 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_520 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_521 = _cvpt_514;   // oc8051_tb.v(104)
    assign _cvpt_523 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_524 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_525 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_526 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_527 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_528 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_529 = _cvpt_522;   // oc8051_tb.v(104)
    assign _cvpt_531 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_532 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_533 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_534 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_535 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_536 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_537 = _cvpt_530;   // oc8051_tb.v(104)
    assign _cvpt_539 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_540 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_541 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_542 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_543 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_544 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_545 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_546 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_547 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_548 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_549 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_550 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_551 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_552 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_553 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_554 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_555 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_556 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_557 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_558 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_559 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_560 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_561 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_562 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_563 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_564 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_565 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_566 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_567 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_568 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_569 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_570 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_571 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_572 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_573 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_574 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_575 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_576 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_577 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_578 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_579 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_580 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_581 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_582 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_583 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_584 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_585 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_586 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_587 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_588 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_589 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_590 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_591 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_592 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_593 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_594 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_595 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_596 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_597 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_598 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_599 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_600 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_601 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_602 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_603 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_604 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_605 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_606 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_607 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_608 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_609 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_610 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_611 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_612 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_613 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_614 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_615 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_616 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_617 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_618 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_619 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_620 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_621 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_622 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_623 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_624 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_625 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_626 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_627 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_628 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_629 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_630 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_631 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_632 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_633 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_634 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_635 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_636 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_637 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_638 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_639 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_640 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_641 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_642 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_643 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_644 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_645 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_646 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_647 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_648 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_649 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_650 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_651 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_652 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_653 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_654 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_655 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_656 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_657 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_658 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_659 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_660 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_661 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_662 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_663 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_664 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_665 = _cvpt_538;   // oc8051_tb.v(104)
    assign _cvpt_666 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_667 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_668 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_669 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_670 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_671 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_672 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_673 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_674 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_675 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_676 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_677 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_678 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_679 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_680 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_681 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_682 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_683 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_684 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_685 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_686 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_687 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_688 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_689 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_690 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_691 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_692 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_693 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_694 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_695 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_696 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_697 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_698 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_699 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_700 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_701 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_702 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_703 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_704 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_705 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_706 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_707 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_708 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_709 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_710 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_711 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_712 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_713 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_714 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_715 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_716 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_717 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_718 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_719 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_720 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_721 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_722 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_723 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_724 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_725 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_726 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_727 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_728 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_729 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_730 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_731 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_732 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_733 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_734 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_735 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_736 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_737 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_738 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_739 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_740 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_741 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_742 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_743 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_744 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_745 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_746 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_747 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_748 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_749 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_750 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_751 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_752 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_753 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_754 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_755 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_756 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_757 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_758 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_759 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_760 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_761 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_762 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_763 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_764 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_765 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_766 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_767 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_768 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_769 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_770 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_771 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_772 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_773 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_774 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_775 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_776 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_777 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_778 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_779 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_780 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_781 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_782 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_783 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_784 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_785 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_786 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_787 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_788 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_789 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_790 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_791 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_792 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_793 = _cvpt_404;   // oc8051_tb.v(104)
    assign _cvpt_795 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_796 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_797 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_798 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_799 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_800 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_801 = _cvpt_794;   // oc8051_tb.v(104)
    assign _cvpt_803 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_804 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_805 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_806 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_807 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_808 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_809 = _cvpt_802;   // oc8051_tb.v(104)
    assign _cvpt_811 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_812 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_813 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_814 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_815 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_816 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_817 = _cvpt_810;   // oc8051_tb.v(104)
    assign _cvpt_819 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_820 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_821 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_822 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_823 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_824 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_825 = _cvpt_818;   // oc8051_tb.v(104)
    assign _cvpt_827 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_828 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_829 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_830 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_831 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_832 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_833 = _cvpt_826;   // oc8051_tb.v(104)
    assign _cvpt_835 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_836 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_837 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_838 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_839 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_840 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_841 = _cvpt_834;   // oc8051_tb.v(104)
    assign _cvpt_843 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_844 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_845 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_846 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_847 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_848 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_849 = _cvpt_842;   // oc8051_tb.v(104)
    assign _cvpt_851 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_852 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_853 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_854 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_855 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_856 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_857 = _cvpt_850;   // oc8051_tb.v(104)
    assign _cvpt_859 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_860 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_861 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_862 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_863 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_864 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_865 = _cvpt_858;   // oc8051_tb.v(104)
    assign _cvpt_867 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_868 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_869 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_870 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_871 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_872 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_873 = _cvpt_866;   // oc8051_tb.v(104)
    assign _cvpt_875 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_876 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_877 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_878 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_879 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_880 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_881 = _cvpt_874;   // oc8051_tb.v(104)
    assign _cvpt_883 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_884 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_885 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_886 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_887 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_888 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_889 = _cvpt_882;   // oc8051_tb.v(104)
    assign _cvpt_891 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_892 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_893 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_894 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_895 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_896 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_897 = _cvpt_890;   // oc8051_tb.v(104)
    assign _cvpt_899 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_900 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_901 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_902 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_903 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_904 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_905 = _cvpt_898;   // oc8051_tb.v(104)
    assign _cvpt_907 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_908 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_909 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_910 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_911 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_912 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_913 = _cvpt_906;   // oc8051_tb.v(104)
    assign _cvpt_915 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_916 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_917 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_918 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_919 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_920 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_921 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_922 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_923 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_924 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_925 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_926 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_927 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_928 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_929 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_930 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_931 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_932 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_933 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_934 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_935 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_936 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_937 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_938 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_939 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_940 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_941 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_942 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_943 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_944 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_945 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_946 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_947 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_948 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_949 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_950 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_951 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_952 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_953 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_954 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_955 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_956 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_957 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_958 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_959 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_960 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_961 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_962 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_963 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_964 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_965 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_966 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_967 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_968 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_969 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_970 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_971 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_972 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_973 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_974 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_975 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_976 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_977 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_978 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_979 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_980 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_981 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_982 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_983 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_984 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_985 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_986 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_987 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_988 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_989 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_990 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_991 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_992 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_993 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_994 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_995 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_996 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_997 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_998 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_999 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1000 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1001 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1002 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1003 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1004 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1005 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1006 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1007 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1008 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1009 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1010 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1011 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1012 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1013 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1014 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1015 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1016 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1017 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1018 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1019 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1020 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1021 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1022 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1023 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1024 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1025 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1026 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1027 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1028 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1029 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1030 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1031 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1032 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1033 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1034 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1035 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1036 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1037 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1038 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1039 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1040 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1041 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1042 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1043 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1044 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1045 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1046 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1047 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1048 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1049 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1050 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1051 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1052 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1053 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1054 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1055 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1056 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1057 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1058 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1059 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1060 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1061 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1062 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1063 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1064 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1065 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1066 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1067 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1068 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1069 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1070 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1071 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1072 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1073 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1074 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1075 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1076 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1077 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1078 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1079 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1080 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1081 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1082 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1083 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1084 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1085 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1086 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1087 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1088 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1089 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1090 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1091 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1092 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1093 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1094 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1095 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1096 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1097 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1098 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1099 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1100 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1101 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1102 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1103 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1104 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1105 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1106 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1107 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1108 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1109 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1110 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1111 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1112 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1113 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1114 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1115 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1116 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1117 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1118 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1119 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1120 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1121 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1122 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1123 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1124 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1125 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1126 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1127 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1128 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1129 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1130 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1131 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1132 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1133 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1134 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1135 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1136 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1137 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1138 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1139 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1140 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1141 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1142 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1143 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1144 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1145 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1146 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1147 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1148 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1149 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1150 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1151 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1152 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1153 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1154 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1155 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1156 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1157 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1158 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1159 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1160 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1161 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1162 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1163 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1164 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1165 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1166 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1167 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1168 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1169 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1170 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1171 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1172 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1173 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1174 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1175 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1176 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1177 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1178 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1179 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1180 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1181 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1182 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1183 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1184 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1185 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1186 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1187 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1188 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1189 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1190 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1191 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1192 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1193 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1194 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1195 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1196 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1197 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1198 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1199 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1200 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1201 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1202 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1203 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1204 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1205 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1206 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1207 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1208 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1210 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1211 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1212 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1213 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1214 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1215 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1216 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1217 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1218 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1219 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1220 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1221 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1222 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1223 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1224 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1225 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1226 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1227 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1228 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1229 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1230 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1231 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1232 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1233 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1234 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1235 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1236 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1237 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1238 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1239 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1240 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1241 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1242 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1243 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1244 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1245 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1246 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_1249 = _cvpt_1247;   // oc8051_tb.v(104)
    assign _cvpt_1250 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1251 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1256 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1257 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1258 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1259 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1260 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1261 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1262 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1263 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1264 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1265 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1266 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1267 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1268 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1269 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1270 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1271 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1272 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1273 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1274 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1275 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1276 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1277 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1278 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1279 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1280 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1281 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1282 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1283 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1284 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1285 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1286 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1287 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1288 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1289 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1290 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1291 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1292 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1293 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1294 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1295 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1296 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1297 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1298 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1299 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1300 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1301 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1302 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1303 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1304 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1305 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1306 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1307 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1308 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1309 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1310 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1311 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1312 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1313 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1314 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1315 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1316 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1317 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1318 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1319 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1320 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1321 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1322 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1323 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1324 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1325 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1326 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1327 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1328 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1329 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1330 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1331 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1332 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1333 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1334 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1335 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1336 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1337 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1338 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1339 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1340 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1341 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1342 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1343 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1344 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1345 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1346 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1347 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1348 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1349 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1350 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1351 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1352 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1353 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1354 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1355 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1356 = _cvpt_1255;   // oc8051_tb.v(104)
    assign _cvpt_1357 = _cvpt_1254;   // oc8051_tb.v(104)
    assign _cvpt_1358 = _cvpt_1253;   // oc8051_tb.v(104)
    assign _cvpt_1359 = _cvpt_1252;   // oc8051_tb.v(104)
    assign _cvpt_1364 = _cvpt_1363;   // oc8051_tb.v(104)
    assign _cvpt_1366 = _cvpt_1365;   // oc8051_tb.v(104)
    assign _cvpt_1368 = _cvpt_1367;   // oc8051_tb.v(104)
    assign _cvpt_1369 = _cvpt_1367;   // oc8051_tb.v(104)
    assign _cvpt_1371 = _cvpt_1370;   // oc8051_tb.v(104)
    assign _cvpt_1372 = _cvpt_1370;   // oc8051_tb.v(104)
    assign _cvpt_1373 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1374 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1375 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1376 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_1379 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1380 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1381 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1382 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1383 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1384 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1385 = _cvpt_1378;   // oc8051_tb.v(104)
    assign _cvpt_1387 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1388 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1389 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1390 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1391 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1392 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1393 = _cvpt_1386;   // oc8051_tb.v(104)
    assign _cvpt_1394 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1395 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1396 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1397 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1398 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1399 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1400 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1402 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1403 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1404 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1405 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1406 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1407 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1408 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1409 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_1410 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_1412 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1413 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1414 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1415 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1416 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1417 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1418 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1419 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1421 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1422 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1423 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1424 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1425 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1426 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1427 = _cvpt_1420;   // oc8051_tb.v(104)
    assign _cvpt_1428 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1429 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1430 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1431 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1432 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1433 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1434 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_1436 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1437 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1438 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1439 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1440 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1441 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1442 = _cvpt_1435;   // oc8051_tb.v(104)
    assign _cvpt_1444 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1445 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1446 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1447 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1448 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1449 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1450 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1452 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1453 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1454 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1455 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1456 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1457 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1458 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1460 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1461 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1462 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1463 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1464 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1465 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1466 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1468 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1469 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1470 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1471 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1472 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1473 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1474 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1476 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1477 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1478 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1479 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1480 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1481 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1482 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1484 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1485 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1486 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1487 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1488 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1489 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1490 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1492 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1493 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1494 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1495 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1496 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1497 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1498 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1500 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1501 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1502 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1503 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1504 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1505 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1506 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1508 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1509 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1510 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1511 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1512 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1513 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1514 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1516 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1517 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1518 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1519 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1520 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1521 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1522 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1524 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1525 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1526 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1527 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1528 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1529 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1530 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1532 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1533 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1534 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1535 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1536 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1537 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1538 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1540 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1541 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1542 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1543 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1544 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1545 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1546 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1548 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1549 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1550 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1551 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1552 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1553 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1554 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1556 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1557 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1558 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1559 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1560 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1561 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1562 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1564 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1565 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1566 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1567 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1568 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1569 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1570 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1572 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1573 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1574 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1575 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1576 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1577 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1578 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1580 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1581 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1582 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1583 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1584 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1585 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1586 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1588 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1589 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1590 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1591 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1592 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1593 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1594 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1596 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1597 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1598 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1599 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1600 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1601 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1602 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1604 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1605 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1606 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1607 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1608 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1609 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1610 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1612 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1613 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1614 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1615 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1616 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1617 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1618 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1620 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1621 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1622 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1623 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1624 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1625 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1626 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1628 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1629 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1630 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1631 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1632 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1633 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1634 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1636 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1637 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1638 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1639 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1640 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1641 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1642 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1644 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1645 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1646 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1647 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1648 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1649 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1650 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1652 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1653 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1654 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1655 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1656 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1657 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1658 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1660 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1661 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1662 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1663 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1664 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1665 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1666 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1668 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1669 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1670 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1671 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1672 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1673 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1674 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1676 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1677 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1678 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1679 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1680 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1681 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1682 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1684 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1685 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1686 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1687 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1688 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1689 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1690 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1692 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1693 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1694 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1695 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1696 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1697 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1698 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1699 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1700 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1701 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1702 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1703 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1704 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1705 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1706 = _cvpt_1443;   // oc8051_tb.v(104)
    assign _cvpt_1707 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1708 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1709 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1710 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1711 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1712 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1713 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1714 = _cvpt_1451;   // oc8051_tb.v(104)
    assign _cvpt_1715 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1716 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1717 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1718 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1719 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1720 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1721 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1722 = _cvpt_1459;   // oc8051_tb.v(104)
    assign _cvpt_1723 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1724 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1725 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1726 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1727 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1728 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1729 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1730 = _cvpt_1467;   // oc8051_tb.v(104)
    assign _cvpt_1731 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1732 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1733 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1734 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1735 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1736 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1737 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1738 = _cvpt_1475;   // oc8051_tb.v(104)
    assign _cvpt_1739 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1740 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1741 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1742 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1743 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1744 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1745 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1746 = _cvpt_1483;   // oc8051_tb.v(104)
    assign _cvpt_1747 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1748 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1749 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1750 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1751 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1752 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1753 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1754 = _cvpt_1491;   // oc8051_tb.v(104)
    assign _cvpt_1755 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1756 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1757 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1758 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1759 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1760 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1761 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1762 = _cvpt_1499;   // oc8051_tb.v(104)
    assign _cvpt_1763 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1764 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1765 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1766 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1767 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1768 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1769 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1770 = _cvpt_1507;   // oc8051_tb.v(104)
    assign _cvpt_1771 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1772 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1773 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1774 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1775 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1776 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1777 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1778 = _cvpt_1515;   // oc8051_tb.v(104)
    assign _cvpt_1779 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1780 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1781 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1782 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1783 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1784 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1785 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1786 = _cvpt_1523;   // oc8051_tb.v(104)
    assign _cvpt_1787 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1788 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1789 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1790 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1791 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1792 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1793 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1794 = _cvpt_1531;   // oc8051_tb.v(104)
    assign _cvpt_1795 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1796 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1797 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1798 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1799 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1800 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1801 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1802 = _cvpt_1539;   // oc8051_tb.v(104)
    assign _cvpt_1803 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1804 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1805 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1806 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1807 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1808 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1809 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1810 = _cvpt_1547;   // oc8051_tb.v(104)
    assign _cvpt_1811 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1812 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1813 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1814 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1815 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1816 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1817 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1818 = _cvpt_1555;   // oc8051_tb.v(104)
    assign _cvpt_1819 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1820 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1821 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1822 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1823 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1824 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1825 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1826 = _cvpt_1563;   // oc8051_tb.v(104)
    assign _cvpt_1827 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1828 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1829 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1830 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1831 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1832 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1833 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1834 = _cvpt_1571;   // oc8051_tb.v(104)
    assign _cvpt_1835 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1836 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1837 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1838 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1839 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1840 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1841 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1842 = _cvpt_1579;   // oc8051_tb.v(104)
    assign _cvpt_1843 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1844 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1845 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1846 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1847 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1848 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1849 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1850 = _cvpt_1587;   // oc8051_tb.v(104)
    assign _cvpt_1851 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1852 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1853 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1854 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1855 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1856 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1857 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1858 = _cvpt_1595;   // oc8051_tb.v(104)
    assign _cvpt_1859 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1860 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1861 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1862 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1863 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1864 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1865 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1866 = _cvpt_1603;   // oc8051_tb.v(104)
    assign _cvpt_1867 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1868 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1869 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1870 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1871 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1872 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1873 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1874 = _cvpt_1611;   // oc8051_tb.v(104)
    assign _cvpt_1875 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1876 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1877 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1878 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1879 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1880 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1881 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1882 = _cvpt_1619;   // oc8051_tb.v(104)
    assign _cvpt_1883 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1884 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1885 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1886 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1887 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1888 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1889 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1890 = _cvpt_1627;   // oc8051_tb.v(104)
    assign _cvpt_1891 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1892 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1893 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1894 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1895 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1896 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1897 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1898 = _cvpt_1635;   // oc8051_tb.v(104)
    assign _cvpt_1899 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1900 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1901 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1902 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1903 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1904 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1905 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1906 = _cvpt_1643;   // oc8051_tb.v(104)
    assign _cvpt_1907 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1908 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1909 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1910 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1911 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1912 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1913 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1914 = _cvpt_1651;   // oc8051_tb.v(104)
    assign _cvpt_1915 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1916 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1917 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1918 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1919 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1920 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1921 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1922 = _cvpt_1659;   // oc8051_tb.v(104)
    assign _cvpt_1923 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1924 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1925 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1926 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1927 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1928 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1929 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1930 = _cvpt_1667;   // oc8051_tb.v(104)
    assign _cvpt_1931 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1932 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1933 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1934 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1935 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1936 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1937 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1938 = _cvpt_1675;   // oc8051_tb.v(104)
    assign _cvpt_1939 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1940 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1941 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1942 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1943 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1944 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1945 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1946 = _cvpt_1683;   // oc8051_tb.v(104)
    assign _cvpt_1947 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1948 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1949 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1950 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1951 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1952 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1953 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1954 = _cvpt_1691;   // oc8051_tb.v(104)
    assign _cvpt_1956 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1957 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1958 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1959 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1960 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1961 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1962 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1963 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1964 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1965 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1966 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1967 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1968 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1969 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1970 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1971 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1972 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1973 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1974 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1975 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1976 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1977 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1978 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1979 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1980 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1981 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1982 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1983 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1984 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1985 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1986 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1987 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1988 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1989 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1990 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1991 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1992 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1993 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1994 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1995 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1996 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1997 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1998 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_1999 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2000 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2001 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2002 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2003 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2004 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2005 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2006 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2007 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2008 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2009 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2010 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2011 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2012 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2013 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2014 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2015 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2016 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2017 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2018 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2019 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2020 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2021 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2022 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2023 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2024 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2025 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2026 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2027 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2028 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2029 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2030 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2031 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2032 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2033 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2034 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2035 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2036 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2037 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2038 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2039 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2040 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2041 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2042 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2043 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2044 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2045 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2046 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2047 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2048 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2049 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2050 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2051 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2052 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2053 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2054 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2055 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2056 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2057 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2058 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2059 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2060 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2061 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2062 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2063 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2064 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2065 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2066 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2067 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2068 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2069 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2070 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2071 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2072 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2073 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2074 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2075 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2076 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2077 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2078 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2079 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2080 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2081 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2082 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2083 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2084 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2085 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2086 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2087 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2088 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2089 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2090 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2091 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2092 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2093 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2094 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2095 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2096 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2097 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2098 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2099 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2100 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2101 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2102 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2103 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2104 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2105 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2106 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2107 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2108 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2109 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2110 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2111 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2112 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2113 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2114 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2115 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2116 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2117 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2118 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2119 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2120 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2121 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2122 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2123 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2124 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2125 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2126 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2127 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2128 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2129 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2130 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2131 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2132 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2133 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2134 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2135 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2136 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2137 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2138 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2139 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2140 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2141 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2142 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2143 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2144 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2145 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2146 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2147 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2148 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2149 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2150 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2151 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2152 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2153 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2154 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2155 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2156 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2157 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2158 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2159 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2160 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2161 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2162 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2163 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2164 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2165 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2166 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2167 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2168 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2169 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2170 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2171 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2172 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2173 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2174 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2175 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2176 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2177 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2178 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2179 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2180 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2181 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2182 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2183 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2184 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2185 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2186 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2187 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2188 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2189 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2190 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2191 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2192 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2193 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2194 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2195 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2196 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2197 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2198 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2199 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2200 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2201 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2202 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2203 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2204 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2205 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2206 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2207 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2208 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2209 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2210 = _cvpt_1955;   // oc8051_tb.v(104)
    assign _cvpt_2212 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2213 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2214 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2215 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2216 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2217 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2218 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2219 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2220 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2221 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2222 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2223 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2224 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2225 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2226 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2227 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2228 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2229 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2230 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2231 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2232 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2233 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2234 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2235 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2236 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2237 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2238 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2239 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2240 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2241 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2242 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2243 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2244 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2245 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2246 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2247 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2248 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2249 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2250 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2251 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2252 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2253 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2254 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2255 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2256 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2257 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2258 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2259 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2260 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2261 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2262 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2263 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2264 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2265 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2266 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2267 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2268 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2269 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2270 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2271 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2272 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2273 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2274 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2275 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2276 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2277 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2278 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2279 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2280 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2281 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2282 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2283 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2284 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2285 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2286 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2287 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2288 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2289 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2290 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2291 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2292 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2293 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2294 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2295 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2296 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2297 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2298 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2299 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2300 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2301 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2302 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2303 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2304 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2305 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2306 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2307 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2308 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2309 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2310 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2311 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2312 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2313 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2314 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2315 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2316 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2317 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2318 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2319 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2320 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2321 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2322 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2323 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2324 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2325 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2326 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2327 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2328 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2329 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2330 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2331 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2332 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2333 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2334 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2335 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2336 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2337 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2338 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2339 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2340 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2341 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2342 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2343 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2344 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2345 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2346 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2347 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2348 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2349 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2350 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2351 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2352 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2353 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2354 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2355 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2356 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2357 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2358 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2359 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2360 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2361 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2362 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2363 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2364 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2365 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2366 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2367 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2368 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2369 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2370 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2371 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2372 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2373 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2374 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2375 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2376 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2377 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2378 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2379 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2380 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2381 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2382 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2383 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2384 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2385 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2386 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2387 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2388 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2389 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2390 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2391 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2392 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2393 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2394 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2395 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2396 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2397 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2398 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2399 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2400 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2401 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2402 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2403 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2404 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2405 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2406 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2407 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2408 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2409 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2410 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2411 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2412 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2413 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2414 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2415 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2416 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2417 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2418 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2419 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2420 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2421 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2422 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2423 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2424 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2425 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2426 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2427 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2428 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2429 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2430 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2431 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2432 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2433 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2434 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2435 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2436 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2437 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2438 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2439 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2440 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2441 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2442 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2443 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2444 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2445 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2446 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2447 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2448 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2449 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2450 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2451 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2452 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2453 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2454 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2455 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2456 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2457 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2458 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2459 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2460 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2461 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2462 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2463 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2464 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2465 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2466 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2467 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2468 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2469 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2470 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2471 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2472 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2473 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2474 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2475 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2476 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2477 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2478 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2479 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2480 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2481 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2482 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2483 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2484 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2485 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2486 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2487 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2488 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2489 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2490 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2491 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2492 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2493 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2494 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2495 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2496 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2497 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2498 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2499 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2500 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2501 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2502 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2503 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2504 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2505 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2506 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2507 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2508 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2509 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2510 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2511 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2512 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2513 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2514 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2515 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2516 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2517 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2518 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2519 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2520 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2521 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2522 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2523 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2524 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2525 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2526 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2527 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2528 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2529 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2530 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2531 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2532 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2533 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2534 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2535 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2536 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2537 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2538 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2539 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2540 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2541 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2542 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2543 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2544 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2545 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2546 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2547 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2548 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2549 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2550 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2551 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2552 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2553 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2554 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2555 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2556 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2557 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2558 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2559 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2560 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2561 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2562 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2563 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2564 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2565 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2566 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2567 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2568 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2569 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2570 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2571 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2572 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2573 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2574 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2575 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2576 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2577 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2578 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2579 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2580 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2581 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2582 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2583 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2584 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2585 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2586 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2587 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2588 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2589 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2590 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2591 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2592 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2593 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2594 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2595 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2596 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2597 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2598 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2599 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2600 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2601 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2602 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2603 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2604 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2605 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2606 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2607 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2608 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2609 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2610 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2611 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2612 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2613 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2614 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2615 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2616 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2617 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2618 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2619 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2620 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2621 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2622 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2623 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2624 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2625 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2626 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2627 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2628 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2629 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2630 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2631 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2632 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2633 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2634 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2635 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2636 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2637 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2638 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2639 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2640 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2641 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2642 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2643 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2644 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2645 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2646 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2647 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2648 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2649 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2650 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2651 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2652 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2653 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2654 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2655 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2656 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2657 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2658 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2659 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2660 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2661 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2662 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2663 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2664 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2665 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2666 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2667 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2668 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2669 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2670 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2671 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2672 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2673 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2674 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2675 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2676 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2677 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2678 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2679 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2680 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2681 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2682 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2683 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2684 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2685 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2686 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2687 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2688 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2689 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2690 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2691 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2692 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2693 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2694 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2695 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2696 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2697 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2698 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2699 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2700 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2701 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2702 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2703 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2704 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2705 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2706 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2707 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2708 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2709 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2710 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2711 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2712 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2713 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2714 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2715 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2716 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2717 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2718 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2719 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2720 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2721 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2722 = _cvpt_2211;   // oc8051_tb.v(104)
    assign _cvpt_2723 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2724 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2725 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2726 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2727 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2728 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2729 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2730 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2731 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2732 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2733 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2734 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2735 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2736 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2737 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2738 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2739 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2740 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2741 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2742 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2743 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2744 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2745 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2746 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2747 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2748 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2749 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2750 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2751 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2752 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2753 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2754 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2755 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2756 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2757 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2758 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2759 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2760 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2761 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2762 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2763 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2764 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2765 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2766 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2767 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2768 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2769 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2770 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2771 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2772 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2773 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2774 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2775 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2776 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2777 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2778 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2779 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2780 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2781 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2782 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2783 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2784 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2785 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2786 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2787 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2788 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2789 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2790 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2791 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2792 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2793 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2794 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2795 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2796 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2797 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2798 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2799 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2800 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2801 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2802 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2803 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2804 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2805 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2806 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2807 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2808 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2809 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2810 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2811 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2812 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2813 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2814 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2815 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2816 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2817 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2818 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2819 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2820 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2821 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2822 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2823 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2824 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2825 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2826 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2827 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2828 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2829 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2830 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2831 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2832 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2833 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2834 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2835 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2836 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2837 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2838 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2839 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2840 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2841 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2842 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2843 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2844 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2845 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2846 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2847 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2848 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2849 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2850 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2851 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2852 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2853 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2854 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2855 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2856 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2857 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2858 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2859 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2860 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2861 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2862 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2863 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2864 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2865 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2866 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2867 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2868 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2869 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2870 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2871 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2872 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2873 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2874 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2875 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2876 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2877 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2878 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2879 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2880 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2881 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2882 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2883 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2884 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2885 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2886 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2887 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2888 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2889 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2890 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2891 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2892 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2893 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2894 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2895 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2896 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2897 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2898 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2899 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2900 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2901 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2902 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2903 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2904 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2905 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2906 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2907 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2908 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2909 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2910 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2911 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2912 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2913 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2914 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2915 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2916 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2917 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2918 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2919 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2920 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2921 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2922 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2923 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2924 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2925 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2926 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2927 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2928 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2929 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2930 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2931 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2932 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2933 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2934 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2935 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2936 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2937 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2938 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2939 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2940 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2941 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2942 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2943 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2944 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2945 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2946 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2947 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2948 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2949 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2950 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2951 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2952 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2953 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2954 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2955 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2956 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2957 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2958 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2959 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2960 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2961 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2962 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2963 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2964 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2965 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2966 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2967 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2968 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2969 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2970 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2971 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2972 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2973 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2974 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2975 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2976 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2977 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2978 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2979 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2980 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2981 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2982 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2983 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2984 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2985 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2986 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2987 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2988 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2989 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2990 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2991 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2992 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2993 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2994 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2995 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2996 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2997 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2998 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_2999 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3000 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3001 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3002 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3003 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3004 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3005 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3006 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3007 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3008 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3009 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3010 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3011 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3012 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3013 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3014 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3015 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3016 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3017 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3018 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3019 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3020 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3021 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3022 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3023 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3024 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3025 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3026 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3027 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3028 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3029 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3030 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3031 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3032 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3033 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3034 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3035 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3036 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3037 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3038 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3039 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3040 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3041 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3042 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3043 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3044 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3045 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3046 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3047 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3048 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3049 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3050 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3051 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3052 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3053 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3054 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3055 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3056 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3057 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3058 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3059 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3060 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3061 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3062 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3063 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3064 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3065 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3066 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3067 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3068 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3069 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3070 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3071 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3072 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3073 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3074 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3075 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3076 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3077 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3078 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3079 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3080 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3081 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3082 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3083 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3084 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3085 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3086 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3087 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3088 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3089 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3090 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3091 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3092 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3093 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3094 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3095 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3096 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3097 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3098 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3099 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3100 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3101 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3102 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3103 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3104 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3105 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3106 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3107 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3108 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3109 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3110 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3111 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3112 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3113 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3114 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3115 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3116 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3117 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3118 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3119 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3120 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3121 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3122 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3123 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3124 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3125 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3126 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3127 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3128 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3129 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3130 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3131 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3132 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3133 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3134 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3135 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3136 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3137 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3138 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3139 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3140 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3141 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3142 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3143 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3144 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3145 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3146 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3147 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3148 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3149 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3150 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3151 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3152 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3153 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3154 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3155 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3156 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3157 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3158 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3159 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3160 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3161 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3162 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3163 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3164 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3165 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3166 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3167 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3168 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3169 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3170 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3171 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3172 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3173 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3174 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3175 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3176 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3177 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3178 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3179 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3180 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3181 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3182 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3183 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3184 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3185 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3186 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3187 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3188 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3189 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3190 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3191 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3192 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3193 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3194 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3195 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3196 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3197 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3198 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3199 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3200 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3201 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3202 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3203 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3204 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3205 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3206 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3207 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3208 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3209 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3210 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3211 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3212 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3213 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3214 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3215 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3216 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3217 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3218 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3219 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3220 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3221 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3222 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3223 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3224 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3225 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3226 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3227 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3228 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3229 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3230 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3231 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3232 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3233 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3234 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3235 = _cvpt_1209;   // oc8051_tb.v(104)
    assign _cvpt_3238 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3239 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3240 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3241 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3242 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3243 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3244 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3245 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3246 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3247 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3248 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3249 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3250 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3251 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3252 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3253 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3254 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3255 = _cvpt_3237;   // oc8051_tb.v(104)
    assign _cvpt_3257 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3258 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3259 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3260 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3261 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3262 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3263 = _cvpt_3256;   // oc8051_tb.v(104)
    assign _cvpt_3265 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3266 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3267 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3268 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3269 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3270 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3271 = _cvpt_3264;   // oc8051_tb.v(104)
    assign _cvpt_3273 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3274 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3275 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3276 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3277 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3278 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3279 = _cvpt_3272;   // oc8051_tb.v(104)
    assign _cvpt_3281 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3282 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3283 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3284 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3285 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3286 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3287 = _cvpt_3280;   // oc8051_tb.v(104)
    assign _cvpt_3289 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3290 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3291 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3292 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3293 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3294 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3295 = _cvpt_3288;   // oc8051_tb.v(104)
    assign _cvpt_3297 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3298 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3299 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3300 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3301 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3302 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3303 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3304 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3305 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3306 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3307 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3308 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3309 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3310 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3311 = _cvpt_3296;   // oc8051_tb.v(104)
    assign _cvpt_3313 = _cvpt_3312;   // oc8051_tb.v(104)
    assign _cvpt_3315 = _cvpt_3314;   // oc8051_tb.v(104)
    assign _cvpt_3316 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3317 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3318 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3319 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3320 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3321 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3322 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3323 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3324 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3325 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3326 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3327 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3328 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3329 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3330 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3331 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3332 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3333 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3334 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3335 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3336 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3337 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3338 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3339 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3340 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3341 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3342 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3343 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3344 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3345 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3346 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3347 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3348 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3349 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3350 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3351 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3352 = _cvpt_914;   // oc8051_tb.v(104)
    assign _cvpt_3465 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3467 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3468 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3469 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3471 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3472 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3473 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3474 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3475 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3476 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3477 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3479 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3480 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3481 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3482 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3483 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3484 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3485 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3486 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3487 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3488 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3489 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3490 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3491 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3492 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3493 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3495 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3496 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3497 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3498 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3499 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3500 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3501 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3502 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3503 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3504 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3505 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3506 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3507 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3508 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3509 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3510 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3511 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3512 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3513 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3514 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3515 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3516 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3517 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3518 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3519 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3520 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3521 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3522 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3523 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3524 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3525 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3526 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3527 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3528 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3529 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3530 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3531 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3532 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3533 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3534 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3535 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3536 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3537 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3538 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3539 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3540 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3541 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3542 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3543 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3544 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3545 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3546 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3547 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3548 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3549 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3550 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3551 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3552 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3553 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3554 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3555 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3556 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3557 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3558 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3559 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3560 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3561 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3562 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3563 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3564 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3565 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3566 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3567 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3568 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3569 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3570 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3571 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3572 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3573 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3574 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3575 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3576 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3577 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3578 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3579 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3580 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3581 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3582 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3583 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3584 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3585 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3586 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3587 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3588 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3589 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3590 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3591 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3592 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3593 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3594 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3595 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3596 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3597 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3598 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3599 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3600 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3601 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3602 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3603 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3604 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3605 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3606 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3607 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3608 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3609 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3610 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3611 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3612 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3613 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3614 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3615 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3616 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3617 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3618 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3619 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3620 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3621 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3622 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3623 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3624 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3625 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3626 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3627 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3628 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3629 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3630 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3631 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3632 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3633 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3634 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3635 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3636 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3637 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3638 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3639 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3640 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3641 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3642 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3643 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3644 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3645 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3646 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3647 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3648 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3649 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3650 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3651 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3652 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3653 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3654 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3655 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3656 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3657 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3658 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3659 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3660 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3661 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3662 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3663 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3664 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3665 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3666 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3667 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3668 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3669 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3670 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3671 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3672 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3673 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3674 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3675 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3676 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3677 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3678 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3679 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3680 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3681 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3682 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3683 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3684 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3685 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3686 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3687 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3688 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3689 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3690 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3691 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3692 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3693 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3694 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3695 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3696 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3697 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3698 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3699 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3700 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3701 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3702 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3703 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3704 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3705 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3707 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3708 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3709 = _cvpt_3706;   // oc8051_tb.v(104)
    assign _cvpt_3711 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3712 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3713 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3714 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3715 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3716 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3717 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3718 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3719 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3720 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3721 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3722 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3723 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3724 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3725 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3726 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3727 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3728 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3729 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3730 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3731 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3732 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3733 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3734 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3735 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3736 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3737 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3738 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3739 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3740 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3741 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3742 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3743 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3744 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3745 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3746 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3747 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3748 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3749 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3750 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3751 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3752 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3753 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3754 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3755 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3756 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3757 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3758 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3759 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3760 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3761 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3762 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3763 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3764 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3765 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3766 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3767 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3768 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3769 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3770 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3771 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3772 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3773 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3774 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3775 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3776 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3777 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3778 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3779 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3780 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3781 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3782 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3783 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3784 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3785 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3786 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3787 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3788 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3789 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3790 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3791 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3792 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3793 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3794 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3795 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3796 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3797 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3798 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3799 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3800 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3801 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3802 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3803 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3804 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3805 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3806 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3807 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3808 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3809 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3810 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3811 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3812 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3813 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3814 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3815 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3816 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3817 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3818 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3819 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3820 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3821 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3822 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3823 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3824 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3825 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3826 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3827 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3828 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3829 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3830 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3831 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3832 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3833 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3834 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3835 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3836 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3837 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3838 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3839 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3840 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3841 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3842 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3843 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3844 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3845 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3846 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3847 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3848 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3849 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3850 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3851 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3852 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3853 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3854 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3855 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3856 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3857 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3858 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3859 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3860 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3861 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3862 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3863 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3864 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3865 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3866 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3867 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3868 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3869 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3870 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3871 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3872 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3873 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3874 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3875 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3876 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3877 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3878 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3879 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3880 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3881 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3882 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3883 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3884 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3885 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3886 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3887 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3888 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3889 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3890 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3891 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3892 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3893 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3894 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3895 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3896 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3897 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3898 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3899 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3900 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3901 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3902 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3903 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3904 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3905 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3906 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3907 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3908 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3909 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3910 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3911 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3912 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3913 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3914 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3915 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3916 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3917 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3918 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3919 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3920 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3921 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3922 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3923 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3924 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3925 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3926 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3927 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3928 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3929 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3930 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3931 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3932 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3933 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3934 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3935 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3936 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3937 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3938 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3939 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3940 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3941 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3942 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3943 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3944 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3945 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3946 = _cvpt_1377;   // oc8051_tb.v(104)
    assign _cvpt_3947 = _cvpt_3466;   // oc8051_tb.v(104)
    assign _cvpt_3948 = _cvpt_3470;   // oc8051_tb.v(104)
    assign _cvpt_3949 = _cvpt_3478;   // oc8051_tb.v(104)
    assign _cvpt_3950 = _cvpt_3494;   // oc8051_tb.v(104)
    assign _cvpt_3951 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3952 = _cvpt_3706;   // oc8051_tb.v(104)
    assign _cvpt_3953 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3954 = _cvpt_1401;   // oc8051_tb.v(104)
    assign _cvpt_3955 = _cvpt_3706;   // oc8051_tb.v(104)
    assign _cvpt_3956 = _cvpt_3710;   // oc8051_tb.v(104)
    assign _cvpt_3957 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3959 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3960 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3961 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3963 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3964 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3965 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3966 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3967 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3968 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3969 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_3971 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3972 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3973 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3974 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3975 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3976 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3977 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_3978 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3979 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3980 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3981 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3982 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3983 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3984 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_3985 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_3987 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3988 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3989 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3990 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3991 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3992 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_3993 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3994 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3995 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3996 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3997 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_3998 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_3999 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4000 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4001 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4002 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4003 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4004 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4005 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4006 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4007 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4008 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4009 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4010 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4011 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4012 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4013 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4014 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4015 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4016 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4017 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4018 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4019 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4020 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4021 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4022 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4023 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4024 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4025 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4026 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4027 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4028 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4029 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4030 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4031 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4032 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4033 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4034 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4035 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4036 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4037 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4038 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4039 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4040 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4041 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4042 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4043 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4044 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4045 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4046 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4047 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4048 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4049 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4050 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4051 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4052 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4053 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4054 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4055 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4056 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4057 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4058 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4059 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4060 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4061 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4062 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4063 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4064 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4065 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4066 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4067 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4068 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4069 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4070 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4071 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4072 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4073 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4074 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4075 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4076 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4077 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4078 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4079 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4080 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4081 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4082 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4083 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4084 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4085 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4086 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4087 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4088 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4089 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4090 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4091 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4092 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4093 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4094 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4095 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4096 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4097 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4098 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4099 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4100 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4101 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4102 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4103 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4104 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4105 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4106 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4107 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4108 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4109 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4110 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4111 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4112 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4113 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4114 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4115 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4116 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4117 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4118 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4119 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4120 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4121 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4122 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4123 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4124 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4125 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4126 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4127 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4128 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4129 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4130 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4131 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4132 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4133 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4134 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4135 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4136 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4137 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4138 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4139 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4140 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4141 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4142 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4143 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4144 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4145 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4146 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4147 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4148 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4149 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4150 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4151 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4152 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4153 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4154 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4155 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4156 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4157 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4158 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4159 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4160 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4161 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4162 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4163 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4164 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4165 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4166 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4167 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4168 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4169 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4170 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4171 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4172 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4173 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4174 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4175 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4176 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4177 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4178 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4179 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4180 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4181 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4182 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4183 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4184 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4185 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4186 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4187 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4188 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4189 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4190 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4191 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4192 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4193 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4194 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4195 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4196 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4197 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4198 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4199 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4200 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4201 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4202 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4203 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4204 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4205 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4206 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4207 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4208 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4209 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4210 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4211 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4212 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4213 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4214 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4215 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4216 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4217 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4218 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4219 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4220 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4221 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4222 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4223 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4224 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4225 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4226 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4227 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4228 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4229 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4230 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4231 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4232 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4233 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4234 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4235 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4236 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4237 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4238 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4239 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4240 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4241 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4242 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4243 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4244 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4245 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4246 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4247 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4248 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4249 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4250 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4251 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4252 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4253 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4254 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4255 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4256 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4257 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4258 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4259 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4260 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4261 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4262 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4263 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4264 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4265 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4266 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4267 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4268 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4269 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4270 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4271 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4272 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4273 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4274 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4275 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4276 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4277 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4278 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4279 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4280 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4281 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4282 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4283 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4284 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4285 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4286 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4287 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4288 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4289 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4290 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4291 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4292 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4293 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4294 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4295 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4296 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4297 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4298 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4299 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4300 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4301 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4302 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4303 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4304 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4305 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4306 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4307 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4308 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4309 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4310 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4311 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4312 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4313 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4314 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4315 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4316 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4317 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4318 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4319 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4320 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4321 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4322 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4323 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4324 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4325 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4326 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4327 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4328 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4329 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4330 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4331 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4332 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4333 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4334 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4335 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4336 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4337 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4338 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4339 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4340 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4341 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4342 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4343 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4344 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4345 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4346 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4347 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4348 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4349 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4350 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4351 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4352 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4353 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4354 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4355 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4356 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4357 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4358 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4359 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4360 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4361 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4362 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4363 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4364 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4365 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4366 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4367 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4368 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4369 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4370 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4371 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4372 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4373 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4374 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4375 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4376 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4377 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4378 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4379 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4380 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4381 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4382 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4383 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4384 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4385 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4386 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4387 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4388 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4389 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4390 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4391 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4392 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4393 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4394 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4395 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4396 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4397 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4398 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4399 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4400 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4401 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4402 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4403 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4404 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4405 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4406 = _cvpt_3986;   // oc8051_tb.v(104)
    assign _cvpt_4407 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4408 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4409 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4410 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4411 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4412 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4413 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4414 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4415 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4416 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4417 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4418 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4419 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4420 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4421 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4422 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4423 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4424 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4425 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4426 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4427 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4428 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4429 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4430 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4431 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4432 = _cvpt_1411;   // oc8051_tb.v(104)
    assign _cvpt_4433 = _cvpt_3958;   // oc8051_tb.v(104)
    assign _cvpt_4434 = _cvpt_3962;   // oc8051_tb.v(104)
    assign _cvpt_4435 = _cvpt_3970;   // oc8051_tb.v(104)
    assign _cvpt_4436 = _cvpt_3986;   // oc8051_tb.v(104)
    assign p3_in[2] = 1'b0;
    assign ea[0] = 1'b1;
    and (\oc8051_top_1/n72 , \oc8051_top_1/wr_o , \oc8051_top_1/n71 ) ;   // oc8051_top.v(503)
    or (\oc8051_top_1/n71 , \oc8051_top_1/n70 , \oc8051_top_1/wr_ind ) ;   // oc8051_top.v(503)
    oc8051_cxrom oc8051_cxrom1 (.clk(clk), .rst(_cvpt_914), .cxrom_addr({cxrom_addr}), 
            .cxrom_data_out({cxrom_data_out}));   // oc8051_tb.v(145)
    oc8051_symbolic_cxrom oc8051_symbolic_cxrom1 (.clk(clk), .rst(_cvpt_914));   // oc8051_tb.v(153)
    not (\oc8051_top_1/n70 , \oc8051_top_1/wr_addr [7]) ;   // oc8051_top.v(503)
    oc8051_ram_top \oc8051_top_1/oc8051_ram_top1  (.clk(clk), .rst(_cvpt_914), 
            .rd_addr({\oc8051_top_1/rd_addr }), .rd_data({\oc8051_top_1/ram_data }), 
            .wr_addr({\oc8051_top_1/wr_addr }), .bit_addr(\oc8051_top_1/bit_addr_o ), 
            .wr_data({\oc8051_top_1/wr_dat }), .wr(\oc8051_top_1/n72 ), 
            .iram({\oc8051_top_1/iram }), .bit_data_in(\oc8051_top_1/desCy ), 
            .bit_data_out(\oc8051_top_1/bit_data ));   // oc8051_top.v(496)
    oc8051_alu \oc8051_top_1/oc8051_alu1  (.rst(_cvpt_914), .clk(clk), .op_code({\oc8051_top_1/alu_op }), 
            .src1({\oc8051_top_1/src1 }), .src2({\oc8051_top_1/src2 }), 
            .src3({\oc8051_top_1/src3 }), .srcCy(\oc8051_top_1/alu_cy ), 
            .srcAc(\oc8051_top_1/srcAc ), .des_acc({\oc8051_top_1/des_acc }), 
            .sub_result({\oc8051_top_1/sub_result }), .des1({\oc8051_top_1/des1 }), 
            .des2({\oc8051_top_1/des2 }), .desCy(\oc8051_top_1/desCy ), 
            .desAc(\oc8051_top_1/desAc ), .desOv(\oc8051_top_1/desOv ), 
            .bit_in(\oc8051_top_1/bit_out ));   // oc8051_top.v(471)
    termination_fsm tfsm0 (.clk(clk), .rst(_cvpt_914), .pout({p0_out}));   // oc8051_tb.v(233)
    termination_fsm tfsm1 (.clk(clk), .rst(_cvpt_914), .pout({p1_out}));   // oc8051_tb.v(244)
    termination_fsm tfsm2 (.clk(clk), .rst(_cvpt_914), .pout({p2_out}));   // oc8051_tb.v(255)
    termination_fsm tfsm3 (.clk(clk), .rst(_cvpt_914), .pout({_cvpt_0, 
            p3_out[6:5], int1, int0, p3_out[2:0]}));   // oc8051_tb.v(266)
    assign \oc8051_xiommu1/proc_data_in [1] = 1'b0;   // oc8051_tb.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(201)
    oc8051_uart_test oc8051_uart_test1 (.clk(clk), .rst(_cvpt_914), .addr({ext_addr[7:0]}), 
            .wr(write_uart), .wr_bit(p3_out[0]), .data_in({data_out}), 
            .data_out({data_out_uart}), .bit_out(p3_in[1]), .rxd(txd), 
            .ow(p3_out[1]), .intr(p3_in[0]), .ack(ack_uart), .stb(stb_o));   // oc8051_tb.v(331)
    and (write_xram, _cvpt_0, write) ;   // oc8051_tb.v(345)
    not (n153, _cvpt_0) ;   // oc8051_tb.v(346)
    and (write_uart, n153, write) ;   // oc8051_tb.v(346)
    assign data_in[7] = _cvpt_0 ? data_out_xram[7] : data_out_uart[7];   // oc8051_tb.v(347)
    assign data_in[6] = _cvpt_0 ? data_out_xram[6] : data_out_uart[6];   // oc8051_tb.v(347)
    assign data_in[5] = _cvpt_0 ? data_out_xram[5] : data_out_uart[5];   // oc8051_tb.v(347)
    assign data_in[4] = _cvpt_0 ? data_out_xram[4] : data_out_uart[4];   // oc8051_tb.v(347)
    assign data_in[3] = _cvpt_0 ? data_out_xram[3] : data_out_uart[3];   // oc8051_tb.v(347)
    assign data_in[2] = _cvpt_0 ? data_out_xram[2] : data_out_uart[2];   // oc8051_tb.v(347)
    assign data_in[1] = _cvpt_0 ? data_out_xram[1] : data_out_uart[1];   // oc8051_tb.v(347)
    assign data_in[0] = _cvpt_0 ? data_out_xram[0] : data_out_uart[0];   // oc8051_tb.v(347)
    assign ack_i = _cvpt_0 ? ack_xram : ack_uart;   // oc8051_tb.v(348)
    oc8051_alu_src_sel \oc8051_top_1/oc8051_alu_src_sel1  (.clk(clk), .rst(_cvpt_914), 
            .rd(\oc8051_top_1/rd ), .sel1({\oc8051_top_1/src_sel1 }), .sel2({\oc8051_top_1/src_sel2 }), 
            .sel3(\oc8051_top_1/src_sel3 ), .acc({\oc8051_top_1/acc }), 
            .ram({\oc8051_top_1/ram_out }), .pc({\oc8051_top_1/pc }), .dptr({\oc8051_top_1/dptr_hi , 
            \oc8051_top_1/dptr_lo }), .op1({\oc8051_top_1/op1_n }), .op2({\oc8051_top_1/op2_n }), 
            .op3({\oc8051_top_1/op3_n }), .src1({\oc8051_top_1/src1 }), 
            .src2({\oc8051_top_1/src2 }), .src3({\oc8051_top_1/src3 }));   // oc8051_top.v(521)
    oc8051_comp \oc8051_top_1/oc8051_comp1  (.sel({\oc8051_top_1/comp_sel }), 
            .eq(\oc8051_top_1/eq ), .b_in(\oc8051_top_1/bit_out ), .cy(\oc8051_top_1/cy ), 
            .acc({\oc8051_top_1/acc }), .des({\oc8051_top_1/sub_result }));   // oc8051_top.v(544)
    oc8051_rom \oc8051_top_1/oc8051_rom1  (.rst(_cvpt_914), .clk(clk), .ea_int(\oc8051_top_1/ea_int ), 
            .cxrom_data_out({cxrom_data_out}), .data_o({\oc8051_top_1/idat_onchip }));   // oc8051_top.v(557)
    oc8051_cy_select \oc8051_top_1/oc8051_cy_select1  (.cy_sel({\oc8051_top_1/cy_sel }), 
            .cy_in(\oc8051_top_1/cy ), .data_in(\oc8051_top_1/bit_out ), 
            .data_out(\oc8051_top_1/alu_cy ));   // oc8051_top.v(582)
    oc8051_indi_addr \oc8051_top_1/oc8051_indi_addr1  (.clk(clk), .rst(_cvpt_914), 
            .wr_addr({\oc8051_top_1/wr_addr }), .data_in({\oc8051_top_1/wr_dat }), 
            .wr(\oc8051_top_1/n72 ), .wr_bit(\oc8051_top_1/bit_addr_o ), 
            .ri_out({\oc8051_top_1/ri }), .sel(\oc8051_top_1/op1_cur [0]), 
            .bank({\oc8051_top_1/bank_sel }), .iram0({\oc8051_top_1/iram [7:0]}), 
            .iram1({\oc8051_top_1/iram [15:8]}), .iram8({\oc8051_top_1/iram [71:64]}), 
            .iram9({\oc8051_top_1/iram [79:72]}));   // oc8051_top.v(588)
    oc8051_memory_interface \oc8051_top_1/oc8051_memory_interface1  (.clk(clk), 
            .rst(_cvpt_914), .wr_i(\oc8051_top_1/wr ), .wr_o(\oc8051_top_1/wr_o ), 
            .wr_bit_i(\oc8051_top_1/bit_addr ), .wr_bit_o(\oc8051_top_1/bit_addr_o ), 
            .wr_dat({\oc8051_top_1/wr_dat }), .des_acc({\oc8051_top_1/des_acc }), 
            .des1({\oc8051_top_1/des1 }), .des2({\oc8051_top_1/des2 }), 
            .rd_addr({\oc8051_top_1/rd_addr }), .wr_addr({\oc8051_top_1/wr_addr }), 
            .wr_ind(\oc8051_top_1/wr_ind ), .bit_in(\oc8051_top_1/bit_data ), 
            .in_ram({\oc8051_top_1/ram_data }), .sfr({\oc8051_top_1/sfr_out }), 
            .sfr_bit(\oc8051_top_1/sfr_bit ), .bit_out(\oc8051_top_1/bit_out ), 
            .iram_out({\oc8051_top_1/ram_out }), .iack_i(\oc8051_top_1/iack_i ), 
            .iadr_o({cxrom_addr}), .idat_i({\oc8051_top_1/idat_i }), .istb_o(\oc8051_top_1/istb_o ), 
            .out_of_rst(\oc8051_top_1/irom_out_of_rst ), .decoder_new_valid_pc(\oc8051_top_1/decoder_new_valid_pc ), 
            .pc_log({\oc8051_top_1/pc_log }), .pc_log_prev({\oc8051_top_1/pc_log_prev }), 
            .idat_onchip({\oc8051_top_1/idat_onchip }), .dadr_o({ext_addr}), 
            .ddat_o({data_out}), .dwe_o(write), .dstb_o(stb_o), .ddat_i({data_in}), 
            .dack_i(ack_i), .rd_sel({\oc8051_top_1/ram_rd_sel }), .wr_sel({\oc8051_top_1/ram_wr_sel }), 
            .rn({\oc8051_top_1/bank_sel , \oc8051_top_1/op1_cur }), .rd_ind(\oc8051_top_1/rd_ind ), 
            .rd(\oc8051_top_1/rd ), .mem_act({\oc8051_top_1/mem_act }), 
            .mem_wait(_cvpt_19), .mem_pc({\oc8051_top_1/mem_pc }), .ea(ea[0]), 
            .ea_int(\oc8051_top_1/ea_int ), .op1_out({\oc8051_top_1/op1_n }), 
            .op2_out({\oc8051_top_1/op2_n }), .op3_out({\oc8051_top_1/op3_n }), 
            .op1({\oc8051_top_1/op1 }), .op2({\oc8051_top_1/op2 }), .op3({\oc8051_top_1/op3 }), 
            .intr(\oc8051_top_1/intr ), .int_v({\oc8051_top_1/int_src }), 
            .int_ack(\oc8051_top_1/int_ack ), .istb(\oc8051_top_1/istb ), 
            .reti(\oc8051_top_1/reti ), .pc_wr_sel({\oc8051_top_1/pc_wr_sel }), 
            .pc_wr(\oc8051_top_1/n76 ), .pc({\oc8051_top_1/pc }), .dpc_ot({dpc_ot}), 
            .sp_w({\oc8051_top_1/sp_w }), .dptr({\oc8051_top_1/dptr_hi , 
            \oc8051_top_1/dptr_lo }), .ri({\oc8051_top_1/ri }), .acc({\oc8051_top_1/acc }), 
            .sp({\oc8051_top_1/sp }), .etr({\oc8051_top_1/etr }));   // oc8051_top.v(609)
    and (\oc8051_top_1/n76 , \oc8051_top_1/pc_wr , \oc8051_top_1/comp_wait ) ;   // oc8051_top.v(682)
    oc8051_sfr \oc8051_top_1/oc8051_sfr1  (.rst(_cvpt_914), .clk(clk), .adr0({\oc8051_top_1/rd_addr }), 
            .adr1({\oc8051_top_1/wr_addr }), .dat0({\oc8051_top_1/sfr_out }), 
            .dat1({\oc8051_top_1/wr_dat }), .dat2({\oc8051_top_1/des2 }), 
            .des_acc({\oc8051_top_1/des_acc }), .we(\oc8051_top_1/n78 ), 
            .bit_in(\oc8051_top_1/desCy ), .bit_out(\oc8051_top_1/sfr_bit ), 
            .wr_bit(\oc8051_top_1/bit_addr_o ), .ram_rd_sel({\oc8051_top_1/ram_rd_sel }), 
            .ram_wr_sel({\oc8051_top_1/ram_wr_sel }), .wr_sfr({\oc8051_top_1/wr_sfr }), 
            .comp_sel({\oc8051_top_1/comp_sel }), .comp_wait(\oc8051_top_1/comp_wait ), 
            .ie({\oc8051_top_1/ie }), .acc({\oc8051_top_1/acc }), .b_reg({\oc8051_top_1/b_reg }), 
            .etr({\oc8051_top_1/etr }), .priv_lvl(priv_lvl), .sp({\oc8051_top_1/sp }), 
            .sp_w({\oc8051_top_1/sp_w }), .bank_sel({\oc8051_top_1/bank_sel }), 
            .desAc(\oc8051_top_1/desAc ), .desOv(\oc8051_top_1/desOv ), 
            .psw_set({\oc8051_top_1/psw_set }), .srcAc(\oc8051_top_1/srcAc ), 
            .cy(\oc8051_top_1/cy ), .psw({\oc8051_top_1/psw }), .p(\oc8051_top_1/p ), 
            .rmw(\oc8051_top_1/rmw ), .p0_out({p0_out}), .p0_in({p0_in}), 
            .p1_out({p1_out}), .p1_in({p1_in}), .p2_out({p2_out}), .p2_in({p2_in}), 
            .p3_out({_cvpt_0, p3_out[6:5], int1, int0, p3_out[2:0]}), 
            .p3_in({p3_in[2], p3_in[2], p3_in[2], p3_in[2], p3_in[2], 
            p3_in[2:0]}), .int_ack(\oc8051_top_1/int_ack ), .intr(\oc8051_top_1/intr ), 
            .int0(int0), .int1(int1), .reti(\oc8051_top_1/reti ), .int_src({\oc8051_top_1/int_src }), 
            .dptr_hi({\oc8051_top_1/dptr_hi }), .dptr_lo({\oc8051_top_1/dptr_lo }), 
            .wait_data(_cvpt_9));   // oc8051_top.v(699)
    not (\oc8051_top_1/n77 , \oc8051_top_1/wr_ind ) ;   // oc8051_top.v(707)
    and (\oc8051_top_1/n78 , \oc8051_top_1/wr_o , \oc8051_top_1/n77 ) ;   // oc8051_top.v(707)
    oc8051_priv_lvl \oc8051_top_1/oc8051_priv_lvl1  (.clk(clk), .rst(_cvpt_914), 
            .enter_su_mode(\oc8051_top_1/enter_su_mode ), .leave_su_mode(\oc8051_top_1/leave_su_mode ), 
            .priv_lvl(priv_lvl), .su_en(ea[0]));   // oc8051_top.v(791)
    not (\oc8051_top_1/oc8051_decoder1/n4 , _cvpt_104) ;   // oc8051_decoder.v(168)
    not (\oc8051_top_1/oc8051_decoder1/n5 , _cvpt_276) ;   // oc8051_decoder.v(168)
    and (\oc8051_top_1/oc8051_decoder1/n6 , \oc8051_top_1/oc8051_decoder1/n4 , 
        \oc8051_top_1/oc8051_decoder1/n5 ) ;   // oc8051_decoder.v(168)
    not (_cvpt_75, _cvpt_9) ;   // oc8051_decoder.v(168)
    and (\oc8051_top_1/rd , \oc8051_top_1/oc8051_decoder1/n6 , _cvpt_75) ;   // oc8051_decoder.v(168)
    and (\oc8051_top_1/istb , \oc8051_top_1/oc8051_decoder1/n5 , \oc8051_top_1/oc8051_decoder1/stb_i ) ;   // oc8051_decoder.v(170)
    assign _cvpt_208 = _cvpt_9 ? 1'b0 : _cvpt_276;   // oc8051_decoder.v(172)
    assign _cvpt_40 = _cvpt_9 ? 1'b0 : _cvpt_104;   // oc8051_decoder.v(172)
    or (\oc8051_top_1/oc8051_decoder1/n13 , _cvpt_104, _cvpt_276) ;   // oc8051_decoder.v(175)
    or (\oc8051_top_1/oc8051_decoder1/n14 , \oc8051_top_1/oc8051_decoder1/n13 , 
        _cvpt_19) ;   // oc8051_decoder.v(175)
    or (_cvpt_11, \oc8051_top_1/oc8051_decoder1/n14 , _cvpt_9) ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n16  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [7] : \oc8051_top_1/op1_n [7];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n17  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [6] : \oc8051_top_1/op1_n [6];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n18  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [5] : \oc8051_top_1/op1_n [5];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n19  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [4] : \oc8051_top_1/op1_n [4];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n20  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [3] : \oc8051_top_1/op1_n [3];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n21  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [2] : \oc8051_top_1/op1_n [2];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n22  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [1] : \oc8051_top_1/op1_n [1];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/oc8051_decoder1/n23  = _cvpt_11 ? \oc8051_top_1/oc8051_decoder1/op [0] : \oc8051_top_1/op1_n [0];   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_d [7] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n16 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_d [6] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n17 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_d [5] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n18 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_d [4] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n19 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_d [3] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n20 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_cur [2] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n21 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_cur [1] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n22 ;   // oc8051_decoder.v(175)
    assign \oc8051_top_1/op1_cur [0] = _cvpt_19 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n23 ;   // oc8051_decoder.v(175)
    not (\oc8051_top_1/oc8051_decoder1/n32 , _cvpt_19) ;   // oc8051_decoder.v(178)
    not (\oc8051_top_1/oc8051_decoder1/n36 , _cvpt_11) ;   // oc8051_decoder.v(178)
    and (\oc8051_top_1/oc8051_decoder1/n37 , \oc8051_top_1/oc8051_decoder1/n32 , 
        \oc8051_top_1/oc8051_decoder1/n36 ) ;   // oc8051_decoder.v(178)
    and (\oc8051_top_1/decoder_new_valid_pc , \oc8051_top_1/oc8051_decoder1/n37 , 
        \oc8051_top_1/irom_out_of_rst ) ;   // oc8051_decoder.v(178)
    assign \oc8051_top_1/alu_op [3] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/alu_op [3];   // oc8051_decoder.v(182)
    assign \oc8051_top_1/alu_op [2] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/alu_op [2];   // oc8051_decoder.v(182)
    assign \oc8051_top_1/alu_op [1] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/alu_op [1];   // oc8051_decoder.v(182)
    assign \oc8051_top_1/alu_op [0] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/alu_op [0];   // oc8051_decoder.v(182)
    assign \oc8051_top_1/wr_sfr [1] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/wr_sfr [1];   // oc8051_decoder.v(183)
    assign \oc8051_top_1/wr_sfr [0] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/wr_sfr [0];   // oc8051_decoder.v(183)
    assign \oc8051_top_1/ram_rd_sel [2] = _cvpt_9 ? \oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [2] : \oc8051_top_1/oc8051_decoder1/ram_rd_sel [2];   // oc8051_decoder.v(184)
    assign \oc8051_top_1/ram_rd_sel [1] = _cvpt_9 ? \oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [1] : \oc8051_top_1/oc8051_decoder1/ram_rd_sel [1];   // oc8051_decoder.v(184)
    assign \oc8051_top_1/ram_rd_sel [0] = _cvpt_9 ? \oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [0] : \oc8051_top_1/oc8051_decoder1/ram_rd_sel [0];   // oc8051_decoder.v(184)
    assign \oc8051_top_1/ram_wr_sel [2] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [2];   // oc8051_decoder.v(185)
    assign \oc8051_top_1/ram_wr_sel [1] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [1];   // oc8051_decoder.v(185)
    assign \oc8051_top_1/ram_wr_sel [0] = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [0];   // oc8051_decoder.v(185)
    assign \oc8051_top_1/wr  = _cvpt_9 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/wr ;   // oc8051_decoder.v(186)
    not (\oc8051_top_1/oc8051_decoder1/n52 , \oc8051_top_1/op1_cur [2]) ;   // oc8051_decoder.v(201)
    not (\oc8051_top_1/oc8051_decoder1/n53 , \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(204)
    not (\oc8051_top_1/oc8051_decoder1/n56 , \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_58/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(210)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(220)
    not (\oc8051_top_1/oc8051_decoder1/n60 , \oc8051_top_1/oc8051_decoder1/n59 ) ;   // oc8051_decoder.v(210)
    not (\oc8051_top_1/oc8051_decoder1/n61 , \oc8051_top_1/eq ) ;   // oc8051_decoder.v(236)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(227)
    not (\oc8051_top_1/oc8051_decoder1/n72 , \oc8051_top_1/op1_d [6]) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(234)
    not (\oc8051_top_1/oc8051_decoder1/n74 , \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(256)
    not (\oc8051_top_1/oc8051_decoder1/n84 , \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_94/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(270)
    not (\oc8051_top_1/oc8051_decoder1/n91 , \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(270)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(284)
    not (\oc8051_top_1/oc8051_decoder1/n102 , \oc8051_top_1/op1_cur [0]) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_116/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(298)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_144/n1 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n83 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_145/n1 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n83 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_147/n1 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n199 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n147 , \oc8051_top_1/oc8051_decoder1/n80 , 
        \oc8051_top_1/oc8051_decoder1/n83 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_148/n1 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/n425 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n1 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_150/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(361)
    and (\oc8051_top_1/oc8051_decoder1/Select_151/n1 , 1'b0, \oc8051_top_1/oc8051_decoder1/n151 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_152/n1 , \oc8051_top_1/oc8051_decoder1/n144 , 
        \oc8051_top_1/oc8051_decoder1/n143 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n1 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(361)
    not (\oc8051_top_1/oc8051_decoder1/n154 , \oc8051_top_1/oc8051_decoder1/n153 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_155/n1 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_156/n1 , \oc8051_top_1/oc8051_decoder1/n83 , 
        \oc8051_top_1/oc8051_decoder1/n80 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_214/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(431)
    not (\oc8051_top_1/oc8051_decoder1/n158 , \oc8051_top_1/oc8051_decoder1/n157 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n159 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/n436 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n208 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n143 ) ;   // oc8051_decoder.v(423)
    or (\oc8051_top_1/oc8051_decoder1/n209 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/n199 ) ;   // oc8051_decoder.v(423)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_216/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(440)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_219/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(449)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_223/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(458)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_227/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(467)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_235/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(485)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_242/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(503)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_247/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(512)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_251/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(521)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_254/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(530)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_257/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(539)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_261/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(548)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_265/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(557)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_269/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(566)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n1 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n1 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n1 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n543 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_549/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n1 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n543 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n1 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/n86 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_552/n1 , \oc8051_top_1/oc8051_decoder1/n446 , 
        _cvpt_41) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n1 , \oc8051_top_1/oc8051_decoder1/n549 , 
        \oc8051_top_1/oc8051_decoder1/n548 ) ;   // oc8051_decoder.v(1223)
    and (\oc8051_top_1/oc8051_decoder1/Select_556/n1 , ea[0], _cvpt_41) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n556 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n436 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_557/n1 , \oc8051_top_1/oc8051_decoder1/n446 , 
        _cvpt_41) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_558/n1 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/n425 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n1 , \oc8051_top_1/oc8051_decoder1/n543 , 
        \oc8051_top_1/oc8051_decoder1/n539 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n1 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/n143 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n1 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/n502 ) ;   // oc8051_decoder.v(1223)
    not (\oc8051_top_1/oc8051_decoder1/n563 , \oc8051_top_1/oc8051_decoder1/n561 ) ;   // oc8051_decoder.v(1223)
    assign \oc8051_top_1/oc8051_decoder1/Mux_565/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n60  : \oc8051_top_1/oc8051_decoder1/n550 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/n565  = _cvpt_41 ? ea[0] : 1'b0;   // oc8051_decoder.v(1223)
    assign \oc8051_top_1/oc8051_decoder1/Mux_566/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n551 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_567/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n552 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_568/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n553 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_569/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n553 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_570/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n557 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_571/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n558 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_572/n1  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_573/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n559 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_574/n1  = _cvpt_40 ? 1'b1 : 1'b1;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_575/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n560 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_576/n1  = _cvpt_40 ? 1'b1 : \oc8051_top_1/oc8051_decoder1/n563 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_577/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n564 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_578/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n565 ;   // oc8051_decoder.v(1225)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_606/n1 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n317 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_610/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_639/n1 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(1411)
    not (\oc8051_top_1/oc8051_decoder1/n612 , \oc8051_top_1/oc8051_decoder1/n611 ) ;   // oc8051_decoder.v(1347)
    not (\oc8051_top_1/oc8051_decoder1/n613 , \oc8051_top_1/oc8051_decoder1/n607 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_640/n1 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_641/n1 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_708/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(1568)
    not (\oc8051_top_1/oc8051_decoder1/n643 , \oc8051_top_1/oc8051_decoder1/n642 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_717/n1 , \oc8051_top_1/oc8051_decoder1/n91 , 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(1590)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n1 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n1 , \oc8051_top_1/oc8051_decoder1/n102 , 
        \oc8051_top_1/oc8051_decoder1/n84 ) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n1 , \oc8051_top_1/op1_cur [0], 
        \oc8051_top_1/op1_cur [1]) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n1 , \oc8051_top_1/oc8051_decoder1/n512 , 
        _cvpt_41) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n1 , \oc8051_top_1/oc8051_decoder1/n543 , 
        \oc8051_top_1/oc8051_decoder1/n1120 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1141/n1 , \oc8051_top_1/oc8051_decoder1/n473 , 
        _cvpt_41) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n1 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n1115 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n1 , \oc8051_top_1/oc8051_decoder1/n1129 , 
        \oc8051_top_1/oc8051_decoder1/n1115 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n1 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1015 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n1 , \oc8051_top_1/oc8051_decoder1/n1129 , 
        \oc8051_top_1/oc8051_decoder1/n539 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n1 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n543 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n1 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1085 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n1 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1115 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n1 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1115 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n1 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/n543 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n1 , \oc8051_top_1/oc8051_decoder1/n1107 , 
        \oc8051_top_1/oc8051_decoder1/n143 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n1 , \oc8051_top_1/oc8051_decoder1/n1107 , 
        \oc8051_top_1/oc8051_decoder1/n1095 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n1 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/n1095 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n1 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n1 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/n1095 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1156/n1 , \oc8051_top_1/oc8051_decoder1/n1115 , 
        \oc8051_top_1/oc8051_decoder1/n1015 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n1 , \oc8051_top_1/oc8051_decoder1/n1129 , 
        \oc8051_top_1/oc8051_decoder1/n539 ) ;   // oc8051_decoder.v(2696)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1158/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n612  : \oc8051_top_1/oc8051_decoder1/n1142 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1159/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n613  : \oc8051_top_1/oc8051_decoder1/n1143 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1160/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n613  : \oc8051_top_1/oc8051_decoder1/n1144 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1161/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1145 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1162/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1146 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1163/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1147 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1164/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n139  : \oc8051_top_1/oc8051_decoder1/n1148 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1165/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n143  : \oc8051_top_1/oc8051_decoder1/n1149 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1166/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n143  : \oc8051_top_1/oc8051_decoder1/n1150 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1167/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n1152 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1168/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1153 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1169/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n456 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1170/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n1140 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1171/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n1141 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1172/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n1151 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1173/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1154 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1174/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1155 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1175/n1  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1156 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1176/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n1157 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1177/n1  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n612  : \oc8051_top_1/oc8051_decoder1/n1158 ;   // oc8051_decoder.v(2698)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1219/n1 , _cvpt_104, _cvpt_276) ;   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1179  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1159  : \oc8051_top_1/src_sel1 [2];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1180  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1160  : \oc8051_top_1/src_sel1 [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1181  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1161  : \oc8051_top_1/src_sel1 [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1182  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1162  : \oc8051_top_1/src_sel2 [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1183  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1163  : \oc8051_top_1/src_sel2 [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1184  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1164  : \oc8051_top_1/oc8051_decoder1/alu_op [3];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1185  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1165  : \oc8051_top_1/oc8051_decoder1/alu_op [2];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1186  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1166  : \oc8051_top_1/oc8051_decoder1/alu_op [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1187  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1167  : \oc8051_top_1/oc8051_decoder1/alu_op [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1188  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1168  : \oc8051_top_1/psw_set [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1189  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1169  : \oc8051_top_1/psw_set [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1190  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1170  : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [2];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1191  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1171  : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1192  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1172  : \oc8051_top_1/oc8051_decoder1/ram_wr_sel [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1193  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1173  : \oc8051_top_1/oc8051_decoder1/wr ;   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1194  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1174  : \oc8051_top_1/cy_sel [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1195  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1175  : \oc8051_top_1/cy_sel [0];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1196  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1176  : \oc8051_top_1/src_sel3 ;   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1197  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1177  : \oc8051_top_1/oc8051_decoder1/wr_sfr [1];   // oc8051_decoder.v(2699)
    assign \oc8051_top_1/oc8051_decoder1/n1198  = _cvpt_75 ? \oc8051_top_1/oc8051_decoder1/n1178  : \oc8051_top_1/oc8051_decoder1/wr_sfr [0];   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1200  (.d(\oc8051_top_1/oc8051_decoder1/n1191 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_wr_sel [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1201  (.d(\oc8051_top_1/oc8051_decoder1/n1192 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_wr_sel [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1202  (.d(\oc8051_top_1/oc8051_decoder1/n1179 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel1 [2]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1203  (.d(\oc8051_top_1/oc8051_decoder1/n1180 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel1 [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1204  (.d(\oc8051_top_1/oc8051_decoder1/n1181 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel1 [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1205  (.d(\oc8051_top_1/oc8051_decoder1/n1182 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel2 [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1206  (.d(\oc8051_top_1/oc8051_decoder1/n1183 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel2 [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1207  (.d(\oc8051_top_1/oc8051_decoder1/n1184 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/alu_op [3]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1208  (.d(\oc8051_top_1/oc8051_decoder1/n1185 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/alu_op [2]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1209  (.d(\oc8051_top_1/oc8051_decoder1/n1186 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/alu_op [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1210  (.d(\oc8051_top_1/oc8051_decoder1/n1187 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/alu_op [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1211  (.d(\oc8051_top_1/oc8051_decoder1/n1193 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/wr ));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1212  (.d(\oc8051_top_1/oc8051_decoder1/n1188 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/psw_set [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1213  (.d(\oc8051_top_1/oc8051_decoder1/n1189 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/psw_set [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1214  (.d(\oc8051_top_1/oc8051_decoder1/n1194 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/cy_sel [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1215  (.d(\oc8051_top_1/oc8051_decoder1/n1195 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/cy_sel [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1216  (.d(\oc8051_top_1/oc8051_decoder1/n1196 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/src_sel3 ));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1217  (.d(\oc8051_top_1/oc8051_decoder1/n1197 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/wr_sfr [1]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1218  (.d(\oc8051_top_1/oc8051_decoder1/n1198 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/wr_sfr [0]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1229  (.d(\oc8051_top_1/oc8051_decoder1/n1221 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [7]));   // oc8051_decoder.v(2707)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2721)
    assign \oc8051_top_1/oc8051_decoder1/n1221  = _cvpt_95 ? \oc8051_top_1/op1_n [7] : \oc8051_top_1/oc8051_decoder1/op [7];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1222  = _cvpt_95 ? \oc8051_top_1/op1_n [6] : \oc8051_top_1/oc8051_decoder1/op [6];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1223  = _cvpt_95 ? \oc8051_top_1/op1_n [5] : \oc8051_top_1/oc8051_decoder1/op [5];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1224  = _cvpt_95 ? \oc8051_top_1/op1_n [4] : \oc8051_top_1/oc8051_decoder1/op [4];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1225  = _cvpt_95 ? \oc8051_top_1/op1_n [3] : \oc8051_top_1/oc8051_decoder1/op [3];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1226  = _cvpt_95 ? \oc8051_top_1/op1_n [2] : \oc8051_top_1/oc8051_decoder1/op [2];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1227  = _cvpt_95 ? \oc8051_top_1/op1_n [1] : \oc8051_top_1/oc8051_decoder1/op [1];   // oc8051_decoder.v(2707)
    assign \oc8051_top_1/oc8051_decoder1/n1228  = _cvpt_95 ? \oc8051_top_1/op1_n [0] : \oc8051_top_1/oc8051_decoder1/op [0];   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1230  (.d(\oc8051_top_1/oc8051_decoder1/n1222 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [6]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1231  (.d(\oc8051_top_1/oc8051_decoder1/n1223 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [5]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1232  (.d(\oc8051_top_1/oc8051_decoder1/n1224 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [4]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1233  (.d(\oc8051_top_1/oc8051_decoder1/n1225 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [3]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1234  (.d(\oc8051_top_1/oc8051_decoder1/n1226 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [2]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1235  (.d(\oc8051_top_1/oc8051_decoder1/n1227 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [1]));   // oc8051_decoder.v(2707)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1236  (.d(\oc8051_top_1/oc8051_decoder1/n1228 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/op [0]));   // oc8051_decoder.v(2707)
    and (_cvpt_106, \oc8051_top_1/oc8051_decoder1/n32 , _cvpt_75) ;   // oc8051_decoder.v(2715)
    not (\oc8051_top_1/oc8051_decoder1/n1241 , \oc8051_top_1/op1_n [0]) ;   // oc8051_decoder.v(2721)
    not (\oc8051_top_1/oc8051_decoder1/n1242 , \oc8051_top_1/op1_n [4]) ;   // oc8051_decoder.v(2721)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2722)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n1 , \oc8051_top_1/oc8051_decoder1/n1246 , 
        \oc8051_top_1/oc8051_decoder1/n1242 ) ;   // oc8051_decoder.v(2723)
    not (\oc8051_top_1/oc8051_decoder1/n1246 , \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2723)
    not (\oc8051_top_1/oc8051_decoder1/n1248 , \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2723)
    not (\oc8051_top_1/oc8051_decoder1/n1249 , \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n1 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2724)
    not (\oc8051_top_1/oc8051_decoder1/n1251 , \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2724)
    not (\oc8051_top_1/oc8051_decoder1/n1252 , \oc8051_top_1/op1_n [2]) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n1 , \oc8051_top_1/oc8051_decoder1/n1246 , 
        \oc8051_top_1/oc8051_decoder1/n1242 ) ;   // oc8051_decoder.v(2728)
    not (\oc8051_top_1/oc8051_decoder1/n1272 , \oc8051_top_1/op1_n [6]) ;   // oc8051_decoder.v(2728)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n1 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n1 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n1 , \oc8051_top_1/oc8051_decoder1/n1241 , 
        \oc8051_top_1/oc8051_decoder1/n1251 ) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n1 , \oc8051_top_1/op1_n [0], 
        \oc8051_top_1/op1_n [1]) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n1 , \oc8051_top_1/oc8051_decoder1/n1354 , 
        \oc8051_top_1/oc8051_decoder1/n1351 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n1 , \oc8051_top_1/oc8051_decoder1/n1348 , 
        \oc8051_top_1/oc8051_decoder1/n1344 ) ;   // oc8051_decoder.v(2752)
    assign \oc8051_top_1/oc8051_decoder1/n1360  = _cvpt_103 ? _cvpt_276 : 1'b1;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1361/n1 , \oc8051_top_1/oc8051_decoder1/n1354 , 
        \oc8051_top_1/oc8051_decoder1/n1324 ) ;   // oc8051_decoder.v(2752)
    and (\oc8051_top_1/oc8051_decoder1/Select_1362/n1 , _cvpt_104, _cvpt_103) ;   // oc8051_decoder.v(2752)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1363/n1  = _cvpt_104 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1360 ;   // oc8051_decoder.v(2754)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1364/n1  = _cvpt_104 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n1363 ;   // oc8051_decoder.v(2754)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n1 , \oc8051_top_1/oc8051_decoder1/n469 , 
        \oc8051_top_1/oc8051_decoder1/n477 ) ;   // oc8051_decoder.v(2785)
    assign \oc8051_top_1/oc8051_decoder1/n1366  = _cvpt_106 ? \oc8051_top_1/oc8051_decoder1/n1364  : _cvpt_276;   // oc8051_decoder.v(2755)
    assign \oc8051_top_1/oc8051_decoder1/n1367  = _cvpt_106 ? \oc8051_top_1/oc8051_decoder1/n1365  : _cvpt_104;   // oc8051_decoder.v(2755)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1369  (.d(\oc8051_top_1/oc8051_decoder1/n1367 ), 
            .clk(clk), .s(_cvpt_914), .r(1'b0), .q(_cvpt_104));   // oc8051_decoder.v(2755)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1371  (.d(\oc8051_top_1/pc [15]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [15]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1372  (.d(\oc8051_top_1/pc [14]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [14]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1373  (.d(\oc8051_top_1/pc [13]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [13]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1374  (.d(\oc8051_top_1/pc [12]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [12]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1375  (.d(\oc8051_top_1/pc [11]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [11]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1376  (.d(\oc8051_top_1/pc [10]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [10]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1377  (.d(\oc8051_top_1/pc [9]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [9]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1378  (.d(\oc8051_top_1/pc [8]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [8]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1379  (.d(\oc8051_top_1/pc [7]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [7]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1380  (.d(\oc8051_top_1/pc [6]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [6]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1381  (.d(\oc8051_top_1/pc [5]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [5]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1382  (.d(\oc8051_top_1/pc [4]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [4]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1383  (.d(\oc8051_top_1/pc [3]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [3]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1384  (.d(\oc8051_top_1/pc [2]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [2]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1385  (.d(\oc8051_top_1/pc [1]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [1]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1386  (.d(\oc8051_top_1/pc [0]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/mem_pc [0]));   // oc8051_decoder.v(2765)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1425  (.d(\oc8051_top_1/oc8051_decoder1/n1422 ), 
            .clk(clk), .s(_cvpt_914), .r(1'b0), .q(\oc8051_top_1/mem_act [2]));   // oc8051_decoder.v(2785)
    not (_cvpt_108, \oc8051_top_1/rd ) ;   // oc8051_decoder.v(2774)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1418/n1 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1419/n1 , \oc8051_top_1/oc8051_decoder1/n317 , 
        \oc8051_top_1/oc8051_decoder1/n323 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1420/n1 , \oc8051_top_1/oc8051_decoder1/n482 , 
        \oc8051_top_1/oc8051_decoder1/n323 ) ;   // oc8051_decoder.v(2785)
    assign \oc8051_top_1/oc8051_decoder1/n1422  = _cvpt_108 ? 1'b1 : \oc8051_top_1/oc8051_decoder1/n1419 ;   // oc8051_decoder.v(2785)
    assign \oc8051_top_1/oc8051_decoder1/n1423  = _cvpt_108 ? 1'b1 : \oc8051_top_1/oc8051_decoder1/n1420 ;   // oc8051_decoder.v(2785)
    assign \oc8051_top_1/oc8051_decoder1/n1424  = _cvpt_108 ? 1'b1 : \oc8051_top_1/oc8051_decoder1/n1421 ;   // oc8051_decoder.v(2785)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1426  (.d(\oc8051_top_1/oc8051_decoder1/n1423 ), 
            .clk(clk), .s(_cvpt_914), .r(1'b0), .q(\oc8051_top_1/mem_act [1]));   // oc8051_decoder.v(2785)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1427  (.d(\oc8051_top_1/oc8051_decoder1/n1424 ), 
            .clk(clk), .s(_cvpt_914), .r(1'b0), .q(\oc8051_top_1/mem_act [0]));   // oc8051_decoder.v(2785)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1429  (.d(\oc8051_top_1/oc8051_decoder1/ram_rd_sel [2]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [2]));   // oc8051_decoder.v(2794)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1430  (.d(\oc8051_top_1/oc8051_decoder1/ram_rd_sel [1]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [1]));   // oc8051_decoder.v(2794)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1431  (.d(\oc8051_top_1/oc8051_decoder1/ram_rd_sel [0]), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_rd_sel_r [0]));   // oc8051_decoder.v(2794)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1199  (.d(\oc8051_top_1/oc8051_decoder1/n1190 ), 
            .clk(clk), .s(1'b0), .r(_cvpt_914), .q(\oc8051_top_1/oc8051_decoder1/ram_wr_sel [2]));   // oc8051_decoder.v(2699)
    VERIFIC_DFFRS \oc8051_top_1/oc8051_decoder1/i1368  (.d(\oc8051_top_1/oc8051_decoder1/n1366 ), 
            .clk(clk), .s(_cvpt_914), .r(1'b0), .q(_cvpt_276));   // oc8051_decoder.v(2755)
    and (_cvpt_151, stb_o, \oc8051_xiommu1/aes_addr_range ) ;   // oc8051_xiommu.v(92)
    and (_cvpt_143, stb_o, \oc8051_xiommu1/sha_addr_range ) ;   // oc8051_xiommu.v(93)
    and (_cvpt_135, stb_o, \oc8051_xiommu1/exp_addr_range ) ;   // oc8051_xiommu.v(94)
    and (_cvpt_127, stb_o, \oc8051_xiommu1/memwr_addr_range ) ;   // oc8051_xiommu.v(95)
    and (_cvpt_119, stb_o, \oc8051_xiommu1/pt_addr_range ) ;   // oc8051_xiommu.v(96)
    and (_cvpt_111, stb_o, \oc8051_xiommu1/ia_addr_range ) ;   // oc8051_xiommu.v(97)
    or (\oc8051_xiommu1/n10 , \oc8051_xiommu1/aes_addr_range , \oc8051_xiommu1/sha_addr_range ) ;   // oc8051_xiommu.v(98)
    or (\oc8051_xiommu1/n11 , \oc8051_xiommu1/n10 , \oc8051_xiommu1/exp_addr_range ) ;   // oc8051_xiommu.v(99)
    or (\oc8051_xiommu1/n12 , \oc8051_xiommu1/n11 , \oc8051_xiommu1/memwr_addr_range ) ;   // oc8051_xiommu.v(99)
    or (\oc8051_xiommu1/n13 , \oc8051_xiommu1/n12 , \oc8051_xiommu1/pt_addr_range ) ;   // oc8051_xiommu.v(100)
    or (\oc8051_xiommu1/n14 , \oc8051_xiommu1/n13 , \oc8051_xiommu1/ia_addr_range ) ;   // oc8051_xiommu.v(100)
    not (\oc8051_xiommu1/n15 , \oc8051_xiommu1/n14 ) ;   // oc8051_xiommu.v(100)
    and (\oc8051_xiommu1/proc1_stb_xram , stb_o, \oc8051_xiommu1/n15 ) ;   // oc8051_xiommu.v(100)
    and (\oc8051_xiommu1/proc0_stb_xram , p3_in[2], \oc8051_xiommu1/n15 ) ;   // oc8051_xiommu.v(103)
    and (\oc8051_xiommu1/write1_xram , \oc8051_xiommu1/proc1_stb_xram , 
        write_xram) ;   // oc8051_xiommu.v(107)
    and (\oc8051_xiommu1/write0_xram , p3_in[2], p3_in[2]) ;   // oc8051_xiommu.v(108)
    and (\oc8051_xiommu1/write_aes , _cvpt_151, write_xram) ;   // oc8051_xiommu.v(109)
    and (\oc8051_xiommu1/write_sha , _cvpt_143, write_xram) ;   // oc8051_xiommu.v(110)
    and (\oc8051_xiommu1/write_exp , _cvpt_135, write_xram) ;   // oc8051_xiommu.v(111)
    and (\oc8051_xiommu1/write_memwr , _cvpt_127, write_xram) ;   // oc8051_xiommu.v(112)
    and (\oc8051_xiommu1/write_pt , _cvpt_119, write_xram) ;   // oc8051_xiommu.v(113)
    or (\oc8051_xiommu1/n31 , \oc8051_xiommu1/proc_ack , \oc8051_xiommu1/ack_aes ) ;   // oc8051_xiommu.v(117)
    or (\oc8051_xiommu1/n32 , \oc8051_xiommu1/n31 , \oc8051_xiommu1/ack_sha ) ;   // oc8051_xiommu.v(117)
    or (\oc8051_xiommu1/n33 , \oc8051_xiommu1/n32 , \oc8051_xiommu1/ack_exp ) ;   // oc8051_xiommu.v(117)
    or (\oc8051_xiommu1/n34 , \oc8051_xiommu1/n33 , \oc8051_xiommu1/ack_memwr ) ;   // oc8051_xiommu.v(117)
    or (\oc8051_xiommu1/n35 , \oc8051_xiommu1/n34 , \oc8051_xiommu1/ack_pt ) ;   // oc8051_xiommu.v(117)
    or (\oc8051_xiommu1/n36 , \oc8051_xiommu1/n35 , \oc8051_xiommu1/ack_ia ) ;   // oc8051_xiommu.v(117)
    and (ack_xram, \oc8051_xiommu1/n36 , _cvpt_1209) ;   // oc8051_xiommu.v(117)
    not (\oc8051_xiommu1/n45 , _cvpt_1209) ;   // oc8051_xiommu.v(118)
    and (\oc8051_xiommu1/proc0_ack , \oc8051_xiommu1/n36 , \oc8051_xiommu1/n45 ) ;   // oc8051_xiommu.v(118)
    assign \oc8051_xiommu1/n47  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [7] : \oc8051_xiommu1/aes_xram_data_in [7];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n48  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [6] : \oc8051_xiommu1/aes_xram_data_in [6];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n49  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [5] : \oc8051_xiommu1/aes_xram_data_in [5];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n50  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [4] : \oc8051_xiommu1/aes_xram_data_in [4];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n51  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [3] : \oc8051_xiommu1/aes_xram_data_in [3];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n52  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [2] : \oc8051_xiommu1/aes_xram_data_in [2];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n53  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [1] : \oc8051_xiommu1/aes_xram_data_in [1];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n54  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [0] : \oc8051_xiommu1/aes_xram_data_in [0];   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n55  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [7] : \oc8051_xiommu1/n47 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n56  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [6] : \oc8051_xiommu1/n48 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n57  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [5] : \oc8051_xiommu1/n49 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n58  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [4] : \oc8051_xiommu1/n50 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n59  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [3] : \oc8051_xiommu1/n51 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n60  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [2] : \oc8051_xiommu1/n52 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n61  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [1] : \oc8051_xiommu1/n53 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n62  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [0] : \oc8051_xiommu1/n54 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n63  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [7] : \oc8051_xiommu1/n55 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n64  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [6] : \oc8051_xiommu1/n56 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n65  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [5] : \oc8051_xiommu1/n57 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n66  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [4] : \oc8051_xiommu1/n58 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n67  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [3] : \oc8051_xiommu1/n59 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n68  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [2] : \oc8051_xiommu1/n60 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n69  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [1] : \oc8051_xiommu1/n61 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n70  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [0] : \oc8051_xiommu1/n62 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n71  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [7] : \oc8051_xiommu1/n63 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n72  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [6] : \oc8051_xiommu1/n64 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n73  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [5] : \oc8051_xiommu1/n65 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n74  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [4] : \oc8051_xiommu1/n66 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n75  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [3] : \oc8051_xiommu1/n67 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n76  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [2] : \oc8051_xiommu1/n68 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n77  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [1] : \oc8051_xiommu1/n69 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n78  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [0] : \oc8051_xiommu1/n70 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n79  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [7] : \oc8051_xiommu1/n71 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n80  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [6] : \oc8051_xiommu1/n72 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n81  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [5] : \oc8051_xiommu1/n73 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n82  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [4] : \oc8051_xiommu1/n74 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n83  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [3] : \oc8051_xiommu1/n75 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n84  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [2] : \oc8051_xiommu1/n76 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n85  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [1] : \oc8051_xiommu1/n77 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n86  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [0] : \oc8051_xiommu1/n78 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[7] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [7] : \oc8051_xiommu1/n79 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[6] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [6] : \oc8051_xiommu1/n80 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[5] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [5] : \oc8051_xiommu1/n81 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[4] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [4] : \oc8051_xiommu1/n82 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[3] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [3] : \oc8051_xiommu1/n83 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[2] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [2] : \oc8051_xiommu1/n84 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[1] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [1] : \oc8051_xiommu1/n85 ;   // oc8051_xiommu.v(137)
    assign data_out_xram[0] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [0] : \oc8051_xiommu1/n86 ;   // oc8051_xiommu.v(137)
    assign \oc8051_xiommu1/n95  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [7] : \oc8051_xiommu1/aes_xram_data_in [7];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n96  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [6] : \oc8051_xiommu1/aes_xram_data_in [6];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n97  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [5] : \oc8051_xiommu1/aes_xram_data_in [5];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n98  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [4] : \oc8051_xiommu1/aes_xram_data_in [4];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n99  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [3] : \oc8051_xiommu1/aes_xram_data_in [3];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n100  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [2] : \oc8051_xiommu1/aes_xram_data_in [2];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n101  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [1] : \oc8051_xiommu1/aes_xram_data_in [1];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n102  = _cvpt_111 ? \oc8051_xiommu1/data_out_ia [0] : \oc8051_xiommu1/aes_xram_data_in [0];   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n103  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [7] : \oc8051_xiommu1/n95 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n104  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [6] : \oc8051_xiommu1/n96 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n105  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [5] : \oc8051_xiommu1/n97 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n106  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [4] : \oc8051_xiommu1/n98 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n107  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [3] : \oc8051_xiommu1/n99 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n108  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [2] : \oc8051_xiommu1/n100 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n109  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [1] : \oc8051_xiommu1/n101 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n110  = _cvpt_119 ? \oc8051_xiommu1/data_out_pt [0] : \oc8051_xiommu1/n102 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n111  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [7] : \oc8051_xiommu1/n103 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n112  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [6] : \oc8051_xiommu1/n104 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n113  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [5] : \oc8051_xiommu1/n105 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n114  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [4] : \oc8051_xiommu1/n106 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n115  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [3] : \oc8051_xiommu1/n107 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n116  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [2] : \oc8051_xiommu1/n108 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n117  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [1] : \oc8051_xiommu1/n109 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n118  = _cvpt_127 ? \oc8051_xiommu1/data_out_memwr [0] : \oc8051_xiommu1/n110 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n119  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [7] : \oc8051_xiommu1/n111 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n120  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [6] : \oc8051_xiommu1/n112 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n121  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [5] : \oc8051_xiommu1/n113 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n122  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [4] : \oc8051_xiommu1/n114 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n123  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [3] : \oc8051_xiommu1/n115 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n124  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [2] : \oc8051_xiommu1/n116 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n125  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [1] : \oc8051_xiommu1/n117 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n126  = _cvpt_135 ? \oc8051_xiommu1/data_out_exp [0] : \oc8051_xiommu1/n118 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n127  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [7] : \oc8051_xiommu1/n119 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n128  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [6] : \oc8051_xiommu1/n120 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n129  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [5] : \oc8051_xiommu1/n121 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n130  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [4] : \oc8051_xiommu1/n122 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n131  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [3] : \oc8051_xiommu1/n123 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n132  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [2] : \oc8051_xiommu1/n124 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n133  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [1] : \oc8051_xiommu1/n125 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/n134  = _cvpt_143 ? \oc8051_xiommu1/data_out_sha [0] : \oc8051_xiommu1/n126 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [7] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [7] : \oc8051_xiommu1/n127 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [6] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [6] : \oc8051_xiommu1/n128 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [5] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [5] : \oc8051_xiommu1/n129 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [4] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [4] : \oc8051_xiommu1/n130 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [3] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [3] : \oc8051_xiommu1/n131 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [2] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [2] : \oc8051_xiommu1/n132 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [1] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [1] : \oc8051_xiommu1/n133 ;   // oc8051_xiommu.v(144)
    assign \oc8051_xiommu1/proc0_data_out [0] = _cvpt_151 ? \oc8051_xiommu1/data_out_aes [0] : \oc8051_xiommu1/n134 ;   // oc8051_xiommu.v(144)
    sha_top \oc8051_xiommu1/sha_top_i  (.clk(clk), .rst(_cvpt_914), .wr(\oc8051_xiommu1/write_sha ), 
            .addr({\oc8051_xiommu1/proc_addr }), .data_in({\oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1:0]}), 
            .data_out({\oc8051_xiommu1/data_out_sha }), .ack(\oc8051_xiommu1/ack_sha ), 
            .stb(_cvpt_143), .in_addr_range(\oc8051_xiommu1/sha_addr_range ), 
            .xram_addr({\oc8051_xiommu1/sha_xram_addr }), .xram_data_out({\oc8051_xiommu1/sha_xram_data_out }), 
            .xram_data_in({\oc8051_xiommu1/aes_xram_data_in }), .xram_ack(\oc8051_xiommu1/sha_xram_ack ), 
            .xram_stb(\oc8051_xiommu1/sha_xram_stb ), .xram_wr(\oc8051_xiommu1/sha_xram_wr ), 
            .sha_state({\oc8051_xiommu1/sha_state }), .sha_rdaddr({\oc8051_xiommu1/sha_rdaddr }), 
            .sha_wraddr({\oc8051_xiommu1/sha_wraddr }), .sha_len({\oc8051_xiommu1/sha_len }), 
            .sha_step(\oc8051_xiommu1/sha_step ), .sha_core_assumps_valid(\oc8051_xiommu1/sha_core_assumps_valid ));   // oc8051_xiommu.v(187)
    modexp_top \oc8051_xiommu1/modexp_top_i  (.clk(clk), .rst(_cvpt_914), 
            .wr(\oc8051_xiommu1/write_exp ), .addr({\oc8051_xiommu1/proc_addr }), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/data_out_exp }), 
            .ack(\oc8051_xiommu1/ack_exp ), .stb(_cvpt_135), .in_addr_range(\oc8051_xiommu1/exp_addr_range ), 
            .xram_addr({\oc8051_xiommu1/exp_xram_addr }), .xram_data_out({\oc8051_xiommu1/exp_xram_data_out }), 
            .xram_data_in({\oc8051_xiommu1/aes_xram_data_in }), .xram_ack(\oc8051_xiommu1/exp_xram_ack ), 
            .xram_stb(\oc8051_xiommu1/exp_xram_stb ), .xram_wr(\oc8051_xiommu1/exp_xram_wr ), 
            .exp_state({\oc8051_xiommu1/exp_state }), .exp_addr({\oc8051_xiommu1/exp_addr }), 
            .exp_step(\oc8051_xiommu1/exp_step ), .exp_m({\oc8051_xiommu1/exp_m }), 
            .exp_exp({\oc8051_xiommu1/exp_exp }), .exp_n({\oc8051_xiommu1/exp_n }), 
            .exp_valid(\oc8051_xiommu1/exp_valid ));   // oc8051_xiommu.v(219)
    mem_wr \oc8051_xiommu1/memwr_i  (.clk(clk), .rst(_cvpt_914), .wr(\oc8051_xiommu1/write_memwr ), 
           .addr({ext_addr}), .data_in({data_out}), .data_out({\oc8051_xiommu1/data_out_memwr }), 
           .ack(\oc8051_xiommu1/ack_memwr ), .stb(_cvpt_127), .in_addr_range(\oc8051_xiommu1/memwr_addr_range ), 
           .xram_addr({\oc8051_xiommu1/memwr_xram_addr }), .xram_data_out({\oc8051_xiommu1/memwr_xram_data_out }), 
           .xram_data_in({\oc8051_xiommu1/aes_xram_data_in }), .xram_ack(\oc8051_xiommu1/memwr_xram_ack ), 
           .xram_stb(\oc8051_xiommu1/memwr_xram_stb ), .xram_wr(\oc8051_xiommu1/memwr_xram_wr ), 
           .memwr_state({\oc8051_xiommu1/memwr_state }), .memwr_rdaddr({\oc8051_xiommu1/memwr_rdaddr }), 
           .memwr_wraddr({\oc8051_xiommu1/memwr_wraddr }), .memwr_len({\oc8051_xiommu1/memwr_len }), 
           .memwr_step(\oc8051_xiommu1/memwr_step ));   // oc8051_xiommu.v(251)
    oc8051_xram \oc8051_xiommu1/oc8051_xram_i  (.clk(clk), .rst(_cvpt_914), 
            .wr(\oc8051_xiommu1/wr_out ), .wr_en(\oc8051_xiommu1/wr_en ), 
            .addr({_cvpt_3494, _cvpt_3478, _cvpt_3470, _cvpt_3466, _cvpt_1377, 
            _cvpt_3710, _cvpt_3706, _cvpt_1401, \oc8051_xiommu1/addr_out [7:5], 
            _cvpt_3986, _cvpt_3970, _cvpt_3962, _cvpt_3958, _cvpt_1411}), 
            .data_in({\oc8051_xiommu1/memarbiter_data_in }), .data_out({\oc8051_xiommu1/aes_xram_data_in }), 
            .ack(\oc8051_xiommu1/ack_in ), .stb(\oc8051_xiommu1/stb_out ), 
            .rd_en(\oc8051_xiommu1/rd_en ));   // oc8051_xiommu.v(359)
    defparam \oc8051_xiommu1/oc8051_xram_i .DELAY = 1;
    xor (_cvpt_3353, 1'b0, \oc8051_xiommu1/proc_addr [0]) ;   // aes_top.v(94)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n2 ) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n5 ) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_53/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n6 ) ;   // oc8051_decoder.v(201)
    not (\oc8051_top_1/oc8051_decoder1/n139 , \oc8051_top_1/oc8051_decoder1/reduce_nor_53/n7 ) ;   // oc8051_decoder.v(201)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n2 ) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n5 ) ;   // oc8051_decoder.v(204)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_57/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n6 ) ;   // oc8051_decoder.v(204)
    not (\oc8051_top_1/oc8051_decoder1/n143 , \oc8051_top_1/oc8051_decoder1/reduce_nor_57/n7 ) ;   // oc8051_decoder.v(204)
    not (\oc8051_top_1/oc8051_decoder1/n59 , \oc8051_top_1/oc8051_decoder1/reduce_nor_58/n1 ) ;   // oc8051_decoder.v(210)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n2 ) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n5 ) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_70/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n6 ) ;   // oc8051_decoder.v(220)
    not (\oc8051_top_1/oc8051_decoder1/n71 , \oc8051_top_1/oc8051_decoder1/reduce_nor_70/n7 ) ;   // oc8051_decoder.v(220)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n2 ) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n5 ) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_72/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n6 ) ;   // oc8051_decoder.v(227)
    not (\oc8051_top_1/oc8051_decoder1/n73 , \oc8051_top_1/oc8051_decoder1/reduce_nor_72/n7 ) ;   // oc8051_decoder.v(227)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n2 ) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n5 ) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_75/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n6 ) ;   // oc8051_decoder.v(234)
    not (\oc8051_top_1/oc8051_decoder1/n76 , \oc8051_top_1/oc8051_decoder1/reduce_nor_75/n7 ) ;   // oc8051_decoder.v(234)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n2 ) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n5 ) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_79/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n6 ) ;   // oc8051_decoder.v(241)
    not (\oc8051_top_1/oc8051_decoder1/n80 , \oc8051_top_1/oc8051_decoder1/reduce_nor_79/n7 ) ;   // oc8051_decoder.v(241)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n2 ) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n5 ) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_82/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n6 ) ;   // oc8051_decoder.v(248)
    not (\oc8051_top_1/oc8051_decoder1/n83 , \oc8051_top_1/oc8051_decoder1/reduce_nor_82/n7 ) ;   // oc8051_decoder.v(248)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n2 ) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n5 ) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_85/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n6 ) ;   // oc8051_decoder.v(256)
    not (\oc8051_top_1/oc8051_decoder1/n86 , \oc8051_top_1/oc8051_decoder1/reduce_nor_85/n7 ) ;   // oc8051_decoder.v(256)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n2 ) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n5 ) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_89/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n6 ) ;   // oc8051_decoder.v(263)
    not (\oc8051_top_1/oc8051_decoder1/n199 , \oc8051_top_1/oc8051_decoder1/reduce_nor_89/n7 ) ;   // oc8051_decoder.v(263)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_94/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(270)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_94/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n2 ) ;   // oc8051_decoder.v(270)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_94/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n3 ) ;   // oc8051_decoder.v(270)
    not (\oc8051_top_1/oc8051_decoder1/n95 , \oc8051_top_1/oc8051_decoder1/reduce_nor_94/n4 ) ;   // oc8051_decoder.v(270)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n1 ) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n4 ) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_100/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n5 ) ;   // oc8051_decoder.v(277)
    not (\oc8051_top_1/oc8051_decoder1/n101 , \oc8051_top_1/oc8051_decoder1/reduce_nor_100/n6 ) ;   // oc8051_decoder.v(277)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n2 ) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n5 ) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_106/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n6 ) ;   // oc8051_decoder.v(284)
    not (\oc8051_top_1/oc8051_decoder1/n107 , \oc8051_top_1/oc8051_decoder1/reduce_nor_106/n7 ) ;   // oc8051_decoder.v(284)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n2 ) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n5 ) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_111/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n6 ) ;   // oc8051_decoder.v(291)
    not (\oc8051_top_1/oc8051_decoder1/n112 , \oc8051_top_1/oc8051_decoder1/reduce_nor_111/n7 ) ;   // oc8051_decoder.v(291)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_116/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(298)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_116/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n2 ) ;   // oc8051_decoder.v(298)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_116/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n3 ) ;   // oc8051_decoder.v(298)
    not (\oc8051_top_1/oc8051_decoder1/n241 , \oc8051_top_1/oc8051_decoder1/reduce_nor_116/n4 ) ;   // oc8051_decoder.v(298)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n2 ) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n5 ) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_122/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n6 ) ;   // oc8051_decoder.v(305)
    not (\oc8051_top_1/oc8051_decoder1/n415 , \oc8051_top_1/oc8051_decoder1/reduce_nor_122/n7 ) ;   // oc8051_decoder.v(305)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n2 ) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n5 ) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_124/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n6 ) ;   // oc8051_decoder.v(312)
    not (\oc8051_top_1/oc8051_decoder1/n425 , \oc8051_top_1/oc8051_decoder1/reduce_nor_124/n7 ) ;   // oc8051_decoder.v(312)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n2 ) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n5 ) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_126/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n6 ) ;   // oc8051_decoder.v(319)
    not (\oc8051_top_1/oc8051_decoder1/n127 , \oc8051_top_1/oc8051_decoder1/reduce_nor_126/n7 ) ;   // oc8051_decoder.v(319)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n2 ) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n5 ) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_132/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n6 ) ;   // oc8051_decoder.v(326)
    not (\oc8051_top_1/oc8051_decoder1/n433 , \oc8051_top_1/oc8051_decoder1/reduce_nor_132/n7 ) ;   // oc8051_decoder.v(326)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n2 ) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n5 ) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_135/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n6 ) ;   // oc8051_decoder.v(333)
    not (\oc8051_top_1/oc8051_decoder1/n436 , \oc8051_top_1/oc8051_decoder1/reduce_nor_135/n7 ) ;   // oc8051_decoder.v(333)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n2 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n433 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n4 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/n425 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n5 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/n112 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n6 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n5 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n6 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n8 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n7 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n9 , \oc8051_top_1/oc8051_decoder1/n107 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n10 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/n86 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n11 , \oc8051_top_1/oc8051_decoder1/n95 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n10 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n12 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n11 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n13 , \oc8051_top_1/oc8051_decoder1/n83 , 
        \oc8051_top_1/oc8051_decoder1/n80 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n14 , \oc8051_top_1/oc8051_decoder1/n73 , 
        \oc8051_top_1/oc8051_decoder1/n71 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n15 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n14 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n16 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n15 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n17 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n16 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_143/n18 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n17 ) ;   // oc8051_decoder.v(361)
    not (\oc8051_top_1/oc8051_decoder1/n144 , \oc8051_top_1/oc8051_decoder1/reduce_nor_143/n18 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_144/n2 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_144/n1 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_144/n3 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/n73 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_144/n4 , \oc8051_top_1/oc8051_decoder1/n80 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_144/n3 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n145 , \oc8051_top_1/oc8051_decoder1/reduce_or_144/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_144/n4 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_145/n2 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_145/n1 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_145/n3 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/n73 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_145/n4 , \oc8051_top_1/oc8051_decoder1/n80 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_145/n3 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n146 , \oc8051_top_1/oc8051_decoder1/reduce_or_145/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_145/n4 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_147/n2 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/n71 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n148 , \oc8051_top_1/oc8051_decoder1/reduce_or_147/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_147/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_148/n2 , \oc8051_top_1/oc8051_decoder1/n83 , 
        \oc8051_top_1/oc8051_decoder1/n73 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n149 , \oc8051_top_1/oc8051_decoder1/reduce_or_148/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_148/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n2 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/n112 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n4 , \oc8051_top_1/oc8051_decoder1/n107 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n5 , \oc8051_top_1/oc8051_decoder1/n80 , 
        \oc8051_top_1/oc8051_decoder1/n76 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n6 , \oc8051_top_1/oc8051_decoder1/n95 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n5 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_149/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n6 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n150 , \oc8051_top_1/oc8051_decoder1/reduce_or_149/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_149/n7 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n151 , \oc8051_top_1/oc8051_decoder1/n144 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_150/n1 ) ;   // oc8051_decoder.v(361)
    and (\oc8051_top_1/oc8051_decoder1/Select_151/n2 , \oc8051_top_1/oc8051_decoder1/n61 , 
        \oc8051_top_1/oc8051_decoder1/n150 ) ;   // oc8051_decoder.v(361)
    and (\oc8051_top_1/oc8051_decoder1/Select_151/n3 , \oc8051_top_1/eq , 
        \oc8051_top_1/oc8051_decoder1/n149 ) ;   // oc8051_decoder.v(361)
    and (\oc8051_top_1/oc8051_decoder1/Select_151/n4 , 1'b1, \oc8051_top_1/oc8051_decoder1/n148 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/Select_151/n5 , \oc8051_top_1/oc8051_decoder1/Select_151/n1 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/Select_151/n6 , \oc8051_top_1/oc8051_decoder1/Select_151/n3 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n4 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n152 , \oc8051_top_1/oc8051_decoder1/Select_151/n5 , 
        \oc8051_top_1/oc8051_decoder1/Select_151/n6 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_152/n2 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/n86 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_152/n3 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_152/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n153 , \oc8051_top_1/oc8051_decoder1/reduce_or_152/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_152/n3 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n2 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n4 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n5 , \oc8051_top_1/oc8051_decoder1/n101 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_154/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n5 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n155 , \oc8051_top_1/oc8051_decoder1/reduce_or_154/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_154/n6 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_155/n2 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/n73 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_155/n3 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_155/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n156 , \oc8051_top_1/oc8051_decoder1/reduce_or_155/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_155/n3 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_156/n2 , \oc8051_top_1/oc8051_decoder1/n76 , 
        \oc8051_top_1/oc8051_decoder1/n73 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/n157 , \oc8051_top_1/oc8051_decoder1/reduce_or_156/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_156/n2 ) ;   // oc8051_decoder.v(361)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_214/n2 , \oc8051_top_1/op1_d [3], 
        \oc8051_top_1/oc8051_decoder1/n74 ) ;   // oc8051_decoder.v(431)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_214/n3 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n2 ) ;   // oc8051_decoder.v(431)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_214/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n3 ) ;   // oc8051_decoder.v(431)
    not (\oc8051_top_1/oc8051_decoder1/n215 , \oc8051_top_1/oc8051_decoder1/reduce_nor_214/n4 ) ;   // oc8051_decoder.v(431)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_216/n2 , \oc8051_top_1/op1_d [3], 
        \oc8051_top_1/op1_d [4]) ;   // oc8051_decoder.v(440)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_216/n3 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n2 ) ;   // oc8051_decoder.v(440)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_216/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n3 ) ;   // oc8051_decoder.v(440)
    not (\oc8051_top_1/oc8051_decoder1/n217 , \oc8051_top_1/oc8051_decoder1/reduce_nor_216/n4 ) ;   // oc8051_decoder.v(440)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_219/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(449)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_219/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n2 ) ;   // oc8051_decoder.v(449)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_219/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n3 ) ;   // oc8051_decoder.v(449)
    not (\oc8051_top_1/oc8051_decoder1/n675 , \oc8051_top_1/oc8051_decoder1/reduce_nor_219/n4 ) ;   // oc8051_decoder.v(449)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_223/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(458)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_223/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n2 ) ;   // oc8051_decoder.v(458)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_223/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n3 ) ;   // oc8051_decoder.v(458)
    not (\oc8051_top_1/oc8051_decoder1/n679 , \oc8051_top_1/oc8051_decoder1/reduce_nor_223/n4 ) ;   // oc8051_decoder.v(458)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_227/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(467)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_227/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n2 ) ;   // oc8051_decoder.v(467)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_227/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n3 ) ;   // oc8051_decoder.v(467)
    not (\oc8051_top_1/oc8051_decoder1/n683 , \oc8051_top_1/oc8051_decoder1/reduce_nor_227/n4 ) ;   // oc8051_decoder.v(467)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_235/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(485)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_235/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n2 ) ;   // oc8051_decoder.v(485)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_235/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n3 ) ;   // oc8051_decoder.v(485)
    not (\oc8051_top_1/oc8051_decoder1/n691 , \oc8051_top_1/oc8051_decoder1/reduce_nor_235/n4 ) ;   // oc8051_decoder.v(485)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_242/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(503)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_242/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n2 ) ;   // oc8051_decoder.v(503)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_242/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n3 ) ;   // oc8051_decoder.v(503)
    not (\oc8051_top_1/oc8051_decoder1/n698 , \oc8051_top_1/oc8051_decoder1/reduce_nor_242/n4 ) ;   // oc8051_decoder.v(503)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_247/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(512)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_247/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n2 ) ;   // oc8051_decoder.v(512)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_247/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n3 ) ;   // oc8051_decoder.v(512)
    not (\oc8051_top_1/oc8051_decoder1/n248 , \oc8051_top_1/oc8051_decoder1/reduce_nor_247/n4 ) ;   // oc8051_decoder.v(512)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_251/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(521)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_251/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n2 ) ;   // oc8051_decoder.v(521)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_251/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n3 ) ;   // oc8051_decoder.v(521)
    not (\oc8051_top_1/oc8051_decoder1/n252 , \oc8051_top_1/oc8051_decoder1/reduce_nor_251/n4 ) ;   // oc8051_decoder.v(521)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_254/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(530)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_254/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n2 ) ;   // oc8051_decoder.v(530)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_254/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n3 ) ;   // oc8051_decoder.v(530)
    not (\oc8051_top_1/oc8051_decoder1/n255 , \oc8051_top_1/oc8051_decoder1/reduce_nor_254/n4 ) ;   // oc8051_decoder.v(530)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_257/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(539)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_257/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n2 ) ;   // oc8051_decoder.v(539)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_257/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n3 ) ;   // oc8051_decoder.v(539)
    not (\oc8051_top_1/oc8051_decoder1/n258 , \oc8051_top_1/oc8051_decoder1/reduce_nor_257/n4 ) ;   // oc8051_decoder.v(539)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_261/n2 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(548)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_261/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n2 ) ;   // oc8051_decoder.v(548)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_261/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n3 ) ;   // oc8051_decoder.v(548)
    not (\oc8051_top_1/oc8051_decoder1/n728 , \oc8051_top_1/oc8051_decoder1/reduce_nor_261/n4 ) ;   // oc8051_decoder.v(548)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_265/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(557)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_265/n3 , \oc8051_top_1/op1_d [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n2 ) ;   // oc8051_decoder.v(557)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_265/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n3 ) ;   // oc8051_decoder.v(557)
    not (\oc8051_top_1/oc8051_decoder1/n732 , \oc8051_top_1/oc8051_decoder1/reduce_nor_265/n4 ) ;   // oc8051_decoder.v(557)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_269/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(566)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_269/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n2 ) ;   // oc8051_decoder.v(566)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_269/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n3 ) ;   // oc8051_decoder.v(566)
    not (\oc8051_top_1/oc8051_decoder1/n270 , \oc8051_top_1/oc8051_decoder1/reduce_nor_269/n4 ) ;   // oc8051_decoder.v(566)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n1 ) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n4 ) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_273/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n5 ) ;   // oc8051_decoder.v(577)
    not (\oc8051_top_1/oc8051_decoder1/n740 , \oc8051_top_1/oc8051_decoder1/reduce_nor_273/n6 ) ;   // oc8051_decoder.v(577)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n1 ) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n4 ) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_278/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n5 ) ;   // oc8051_decoder.v(586)
    not (\oc8051_top_1/oc8051_decoder1/n745 , \oc8051_top_1/oc8051_decoder1/reduce_nor_278/n6 ) ;   // oc8051_decoder.v(586)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n1 ) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n4 ) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_283/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n5 ) ;   // oc8051_decoder.v(595)
    not (\oc8051_top_1/oc8051_decoder1/n750 , \oc8051_top_1/oc8051_decoder1/reduce_nor_283/n6 ) ;   // oc8051_decoder.v(595)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n1 ) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n4 ) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_293/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n5 ) ;   // oc8051_decoder.v(613)
    not (\oc8051_top_1/oc8051_decoder1/n760 , \oc8051_top_1/oc8051_decoder1/reduce_nor_293/n6 ) ;   // oc8051_decoder.v(613)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n1 ) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n4 ) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_296/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n5 ) ;   // oc8051_decoder.v(622)
    not (\oc8051_top_1/oc8051_decoder1/n763 , \oc8051_top_1/oc8051_decoder1/reduce_nor_296/n6 ) ;   // oc8051_decoder.v(622)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n1 ) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n4 ) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_302/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n5 ) ;   // oc8051_decoder.v(631)
    not (\oc8051_top_1/oc8051_decoder1/n303 , \oc8051_top_1/oc8051_decoder1/reduce_nor_302/n6 ) ;   // oc8051_decoder.v(631)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n1 ) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n4 ) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_306/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n5 ) ;   // oc8051_decoder.v(640)
    not (\oc8051_top_1/oc8051_decoder1/n307 , \oc8051_top_1/oc8051_decoder1/reduce_nor_306/n6 ) ;   // oc8051_decoder.v(640)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n1 ) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n4 ) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_311/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n5 ) ;   // oc8051_decoder.v(649)
    not (\oc8051_top_1/oc8051_decoder1/n312 , \oc8051_top_1/oc8051_decoder1/reduce_nor_311/n6 ) ;   // oc8051_decoder.v(649)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n1 ) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n4 ) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_316/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n5 ) ;   // oc8051_decoder.v(658)
    not (\oc8051_top_1/oc8051_decoder1/n317 , \oc8051_top_1/oc8051_decoder1/reduce_nor_316/n6 ) ;   // oc8051_decoder.v(658)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n1 ) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n4 ) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_322/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n5 ) ;   // oc8051_decoder.v(667)
    not (\oc8051_top_1/oc8051_decoder1/n323 , \oc8051_top_1/oc8051_decoder1/reduce_nor_322/n6 ) ;   // oc8051_decoder.v(667)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n1 ) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n4 ) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_326/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n5 ) ;   // oc8051_decoder.v(676)
    not (\oc8051_top_1/oc8051_decoder1/n327 , \oc8051_top_1/oc8051_decoder1/reduce_nor_326/n6 ) ;   // oc8051_decoder.v(676)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n1 ) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n4 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n4 ) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_331/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n5 ) ;   // oc8051_decoder.v(685)
    not (\oc8051_top_1/oc8051_decoder1/n811 , \oc8051_top_1/oc8051_decoder1/reduce_nor_331/n6 ) ;   // oc8051_decoder.v(685)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n1 ) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n4 ) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_336/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n5 ) ;   // oc8051_decoder.v(694)
    not (\oc8051_top_1/oc8051_decoder1/n816 , \oc8051_top_1/oc8051_decoder1/reduce_nor_336/n6 ) ;   // oc8051_decoder.v(694)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n1 ) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n4 ) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_342/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n5 ) ;   // oc8051_decoder.v(703)
    not (\oc8051_top_1/oc8051_decoder1/n822 , \oc8051_top_1/oc8051_decoder1/reduce_nor_342/n6 ) ;   // oc8051_decoder.v(703)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n1 ) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n3 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n4 ) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_347/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n5 ) ;   // oc8051_decoder.v(712)
    not (\oc8051_top_1/oc8051_decoder1/n348 , \oc8051_top_1/oc8051_decoder1/reduce_nor_347/n6 ) ;   // oc8051_decoder.v(712)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n2 ) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n5 ) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_351/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n6 ) ;   // oc8051_decoder.v(723)
    not (\oc8051_top_1/oc8051_decoder1/n831 , \oc8051_top_1/oc8051_decoder1/reduce_nor_351/n7 ) ;   // oc8051_decoder.v(723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n2 ) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n5 ) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_356/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n6 ) ;   // oc8051_decoder.v(732)
    not (\oc8051_top_1/oc8051_decoder1/n839 , \oc8051_top_1/oc8051_decoder1/reduce_nor_356/n7 ) ;   // oc8051_decoder.v(732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n2 ) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n5 ) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_361/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n6 ) ;   // oc8051_decoder.v(741)
    not (\oc8051_top_1/oc8051_decoder1/n848 , \oc8051_top_1/oc8051_decoder1/reduce_nor_361/n7 ) ;   // oc8051_decoder.v(741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n2 ) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n5 ) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_365/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n6 ) ;   // oc8051_decoder.v(750)
    not (\oc8051_top_1/oc8051_decoder1/n852 , \oc8051_top_1/oc8051_decoder1/reduce_nor_365/n7 ) ;   // oc8051_decoder.v(750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n2 ) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n5 ) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_369/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n6 ) ;   // oc8051_decoder.v(759)
    not (\oc8051_top_1/oc8051_decoder1/n856 , \oc8051_top_1/oc8051_decoder1/reduce_nor_369/n7 ) ;   // oc8051_decoder.v(759)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n2 ) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n5 ) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_374/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n6 ) ;   // oc8051_decoder.v(768)
    not (\oc8051_top_1/oc8051_decoder1/n861 , \oc8051_top_1/oc8051_decoder1/reduce_nor_374/n7 ) ;   // oc8051_decoder.v(768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n2 ) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n5 ) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_377/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n6 ) ;   // oc8051_decoder.v(777)
    not (\oc8051_top_1/oc8051_decoder1/n378 , \oc8051_top_1/oc8051_decoder1/reduce_nor_377/n7 ) ;   // oc8051_decoder.v(777)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n2 ) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n5 ) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_381/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n6 ) ;   // oc8051_decoder.v(786)
    not (\oc8051_top_1/oc8051_decoder1/n382 , \oc8051_top_1/oc8051_decoder1/reduce_nor_381/n7 ) ;   // oc8051_decoder.v(786)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n2 ) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n5 ) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_396/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n6 ) ;   // oc8051_decoder.v(813)
    not (\oc8051_top_1/oc8051_decoder1/n397 , \oc8051_top_1/oc8051_decoder1/reduce_nor_396/n7 ) ;   // oc8051_decoder.v(813)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n2 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n5 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_401/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n6 ) ;   // oc8051_decoder.v(822)
    not (\oc8051_top_1/oc8051_decoder1/n402 , \oc8051_top_1/oc8051_decoder1/reduce_nor_401/n7 ) ;   // oc8051_decoder.v(822)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n2 ) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n5 ) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_405/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n6 ) ;   // oc8051_decoder.v(831)
    not (\oc8051_top_1/oc8051_decoder1/n922 , \oc8051_top_1/oc8051_decoder1/reduce_nor_405/n7 ) ;   // oc8051_decoder.v(831)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n2 ) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n5 ) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_417/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n6 ) ;   // oc8051_decoder.v(858)
    not (\oc8051_top_1/oc8051_decoder1/n936 , \oc8051_top_1/oc8051_decoder1/reduce_nor_417/n7 ) ;   // oc8051_decoder.v(858)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n2 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n5 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_422/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n6 ) ;   // oc8051_decoder.v(867)
    not (\oc8051_top_1/oc8051_decoder1/n941 , \oc8051_top_1/oc8051_decoder1/reduce_nor_422/n7 ) ;   // oc8051_decoder.v(867)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n2 ) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n5 ) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_438/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n6 ) ;   // oc8051_decoder.v(949)
    not (\oc8051_top_1/oc8051_decoder1/n439 , \oc8051_top_1/oc8051_decoder1/reduce_nor_438/n7 ) ;   // oc8051_decoder.v(949)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n2 ) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n5 ) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_443/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n6 ) ;   // oc8051_decoder.v(959)
    not (_cvpt_41, \oc8051_top_1/oc8051_decoder1/reduce_nor_443/n7 ) ;   // oc8051_decoder.v(959)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n2 ) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n5 ) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_445/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n6 ) ;   // oc8051_decoder.v(980)
    not (\oc8051_top_1/oc8051_decoder1/n446 , \oc8051_top_1/oc8051_decoder1/reduce_nor_445/n7 ) ;   // oc8051_decoder.v(980)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n2 ) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n5 ) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_451/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n6 ) ;   // oc8051_decoder.v(989)
    not (\oc8051_top_1/oc8051_decoder1/n452 , \oc8051_top_1/oc8051_decoder1/reduce_nor_451/n7 ) ;   // oc8051_decoder.v(989)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n2 ) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n5 ) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_455/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n6 ) ;   // oc8051_decoder.v(998)
    not (\oc8051_top_1/oc8051_decoder1/n456 , \oc8051_top_1/oc8051_decoder1/reduce_nor_455/n7 ) ;   // oc8051_decoder.v(998)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n2 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n5 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_459/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n6 ) ;   // oc8051_decoder.v(1007)
    not (\oc8051_top_1/oc8051_decoder1/n460 , \oc8051_top_1/oc8051_decoder1/reduce_nor_459/n7 ) ;   // oc8051_decoder.v(1007)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n2 ) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n5 ) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_463/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n6 ) ;   // oc8051_decoder.v(1016)
    not (\oc8051_top_1/oc8051_decoder1/n464 , \oc8051_top_1/oc8051_decoder1/reduce_nor_463/n7 ) ;   // oc8051_decoder.v(1016)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n2 ) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n5 ) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_468/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n6 ) ;   // oc8051_decoder.v(1025)
    not (\oc8051_top_1/oc8051_decoder1/n469 , \oc8051_top_1/oc8051_decoder1/reduce_nor_468/n7 ) ;   // oc8051_decoder.v(1025)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n2 ) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n5 ) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_472/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n6 ) ;   // oc8051_decoder.v(1034)
    not (\oc8051_top_1/oc8051_decoder1/n473 , \oc8051_top_1/oc8051_decoder1/reduce_nor_472/n7 ) ;   // oc8051_decoder.v(1034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n2 ) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n5 ) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_476/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n6 ) ;   // oc8051_decoder.v(1043)
    not (\oc8051_top_1/oc8051_decoder1/n477 , \oc8051_top_1/oc8051_decoder1/reduce_nor_476/n7 ) ;   // oc8051_decoder.v(1043)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n2 ) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n5 ) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_481/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n6 ) ;   // oc8051_decoder.v(1052)
    not (\oc8051_top_1/oc8051_decoder1/n482 , \oc8051_top_1/oc8051_decoder1/reduce_nor_481/n7 ) ;   // oc8051_decoder.v(1052)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n2 ) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n5 ) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_489/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n6 ) ;   // oc8051_decoder.v(1070)
    not (\oc8051_top_1/oc8051_decoder1/n490 , \oc8051_top_1/oc8051_decoder1/reduce_nor_489/n7 ) ;   // oc8051_decoder.v(1070)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n2 ) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n5 ) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_492/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n6 ) ;   // oc8051_decoder.v(1079)
    not (\oc8051_top_1/oc8051_decoder1/n493 , \oc8051_top_1/oc8051_decoder1/reduce_nor_492/n7 ) ;   // oc8051_decoder.v(1079)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n2 ) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n5 ) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_496/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n6 ) ;   // oc8051_decoder.v(1088)
    not (\oc8051_top_1/oc8051_decoder1/n497 , \oc8051_top_1/oc8051_decoder1/reduce_nor_496/n7 ) ;   // oc8051_decoder.v(1088)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n2 ) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n5 ) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_501/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n6 ) ;   // oc8051_decoder.v(1097)
    not (\oc8051_top_1/oc8051_decoder1/n502 , \oc8051_top_1/oc8051_decoder1/reduce_nor_501/n7 ) ;   // oc8051_decoder.v(1097)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n2 ) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n5 ) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_504/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n6 ) ;   // oc8051_decoder.v(1106)
    not (\oc8051_top_1/oc8051_decoder1/n505 , \oc8051_top_1/oc8051_decoder1/reduce_nor_504/n7 ) ;   // oc8051_decoder.v(1106)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n2 ) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n5 ) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_508/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n6 ) ;   // oc8051_decoder.v(1115)
    not (\oc8051_top_1/oc8051_decoder1/n509 , \oc8051_top_1/oc8051_decoder1/reduce_nor_508/n7 ) ;   // oc8051_decoder.v(1115)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n2 ) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n5 ) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_511/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n6 ) ;   // oc8051_decoder.v(1124)
    not (\oc8051_top_1/oc8051_decoder1/n512 , \oc8051_top_1/oc8051_decoder1/reduce_nor_511/n7 ) ;   // oc8051_decoder.v(1124)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n2 ) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n5 ) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_523/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n6 ) ;   // oc8051_decoder.v(1151)
    not (\oc8051_top_1/oc8051_decoder1/n524 , \oc8051_top_1/oc8051_decoder1/reduce_nor_523/n7 ) ;   // oc8051_decoder.v(1151)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n2 ) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n5 ) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_528/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n6 ) ;   // oc8051_decoder.v(1169)
    not (\oc8051_top_1/oc8051_decoder1/n1107 , \oc8051_top_1/oc8051_decoder1/reduce_nor_528/n7 ) ;   // oc8051_decoder.v(1169)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n2 ) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n5 ) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_533/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n6 ) ;   // oc8051_decoder.v(1178)
    not (\oc8051_top_1/oc8051_decoder1/n1120 , \oc8051_top_1/oc8051_decoder1/reduce_nor_533/n7 ) ;   // oc8051_decoder.v(1178)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n2 ) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n5 ) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_538/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n6 ) ;   // oc8051_decoder.v(1187)
    not (\oc8051_top_1/oc8051_decoder1/n539 , \oc8051_top_1/oc8051_decoder1/reduce_nor_538/n7 ) ;   // oc8051_decoder.v(1187)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n2 ) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n5 ) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_542/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n6 ) ;   // oc8051_decoder.v(1196)
    not (\oc8051_top_1/oc8051_decoder1/n543 , \oc8051_top_1/oc8051_decoder1/reduce_nor_542/n7 ) ;   // oc8051_decoder.v(1196)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n2 ) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n5 ) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_547/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n6 ) ;   // oc8051_decoder.v(1205)
    not (\oc8051_top_1/oc8051_decoder1/n548 , \oc8051_top_1/oc8051_decoder1/reduce_nor_547/n7 ) ;   // oc8051_decoder.v(1205)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n3 , \oc8051_top_1/oc8051_decoder1/n539 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n5 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/n199 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n6 , \oc8051_top_1/oc8051_decoder1/n512 , 
        \oc8051_top_1/oc8051_decoder1/n509 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n7 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n8 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n7 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n9 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n8 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n10 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/n502 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n11 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n490 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n12 , \oc8051_top_1/oc8051_decoder1/n497 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n11 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n13 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n12 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n14 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n482 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n15 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n16 , \oc8051_top_1/oc8051_decoder1/n477 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n15 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n17 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n16 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n18 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n17 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n19 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n18 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n20 , \oc8051_top_1/oc8051_decoder1/n464 , 
        \oc8051_top_1/oc8051_decoder1/n460 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n21 , \oc8051_top_1/oc8051_decoder1/n452 , 
        \oc8051_top_1/oc8051_decoder1/n446 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n22 , \oc8051_top_1/oc8051_decoder1/n456 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n21 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n23 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n22 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n24 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/n439 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n25 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n26 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n25 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n27 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n26 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n28 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n27 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n29 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n941 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n30 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n31 , \oc8051_top_1/oc8051_decoder1/n936 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n30 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n32 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n31 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n33 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n402 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n34 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n35 , \oc8051_top_1/oc8051_decoder1/n397 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n34 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n36 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n33 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n35 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n37 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n36 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n38 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n37 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n39 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n38 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n40 , \oc8051_top_1/oc8051_decoder1/n382 , 
        \oc8051_top_1/oc8051_decoder1/n378 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n41 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n42 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n41 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n43 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n40 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n42 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n44 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n839 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n45 , \oc8051_top_1/oc8051_decoder1/n348 , 
        \oc8051_top_1/oc8051_decoder1/n822 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n46 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n45 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n47 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n44 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n46 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n48 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n43 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n47 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n49 , \oc8051_top_1/oc8051_decoder1/n816 , 
        \oc8051_top_1/oc8051_decoder1/n811 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n50 , \oc8051_top_1/oc8051_decoder1/n323 , 
        \oc8051_top_1/oc8051_decoder1/n317 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n51 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n50 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n52 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n49 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n51 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n53 , \oc8051_top_1/oc8051_decoder1/n312 , 
        \oc8051_top_1/oc8051_decoder1/n307 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n54 , \oc8051_top_1/oc8051_decoder1/n763 , 
        \oc8051_top_1/oc8051_decoder1/n760 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n55 , \oc8051_top_1/oc8051_decoder1/n303 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n54 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n56 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n53 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n55 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n57 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n52 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n56 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n58 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n48 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n57 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n59 , \oc8051_top_1/oc8051_decoder1/n101 , 
        \oc8051_top_1/oc8051_decoder1/n750 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n60 , \oc8051_top_1/oc8051_decoder1/n740 , 
        \oc8051_top_1/oc8051_decoder1/n270 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n61 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n60 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n62 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n59 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n61 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n63 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n64 , \oc8051_top_1/oc8051_decoder1/n255 , 
        \oc8051_top_1/oc8051_decoder1/n252 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n65 , \oc8051_top_1/oc8051_decoder1/n258 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n64 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n66 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n63 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n65 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n67 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n62 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n66 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n68 , \oc8051_top_1/oc8051_decoder1/n248 , 
        \oc8051_top_1/oc8051_decoder1/n698 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n69 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n70 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n69 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n71 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n68 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n70 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n72 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/n679 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n73 , \oc8051_top_1/oc8051_decoder1/n217 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n74 , \oc8051_top_1/oc8051_decoder1/n675 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n73 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n75 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n72 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n74 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n76 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n71 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n75 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n77 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n67 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n76 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n78 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n58 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n77 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_548/n79 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n39 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n78 ) ;   // oc8051_decoder.v(1223)
    not (\oc8051_top_1/oc8051_decoder1/n549 , \oc8051_top_1/oc8051_decoder1/reduce_nor_548/n79 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_549/n2 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_549/n3 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_549/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n550 , \oc8051_top_1/oc8051_decoder1/reduce_or_549/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_549/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n2 , \oc8051_top_1/oc8051_decoder1/n539 , 
        \oc8051_top_1/oc8051_decoder1/n1120 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n4 , \oc8051_top_1/oc8051_decoder1/n1107 , 
        \oc8051_top_1/oc8051_decoder1/n524 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n5 , \oc8051_top_1/oc8051_decoder1/n86 , 
        \oc8051_top_1/oc8051_decoder1/n512 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n6 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n5 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n7 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n9 , \oc8051_top_1/oc8051_decoder1/n509 , 
        \oc8051_top_1/oc8051_decoder1/n505 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n10 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/n497 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n10 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n12 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n490 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n13 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n456 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n14 , \oc8051_top_1/oc8051_decoder1/n464 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n13 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n14 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n15 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n16 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n18 , \oc8051_top_1/oc8051_decoder1/n452 , 
        \oc8051_top_1/oc8051_decoder1/n436 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n19 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/n425 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n19 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n21 , \oc8051_top_1/oc8051_decoder1/n936 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n22 , \oc8051_top_1/oc8051_decoder1/n402 , 
        \oc8051_top_1/oc8051_decoder1/n397 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n23 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n22 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n23 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n24 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n26 , \oc8051_top_1/oc8051_decoder1/n107 , 
        \oc8051_top_1/oc8051_decoder1/n382 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n27 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n28 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n27 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n28 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n30 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n839 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n31 , \oc8051_top_1/oc8051_decoder1/n312 , 
        \oc8051_top_1/oc8051_decoder1/n252 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n32 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n31 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n32 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n29 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n33 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_550/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n34 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n551 , \oc8051_top_1/oc8051_decoder1/reduce_or_550/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_550/n35 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n2 , \oc8051_top_1/oc8051_decoder1/n509 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n4 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n941 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n5 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n6 , \oc8051_top_1/oc8051_decoder1/n348 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n5 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n7 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n9 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n327 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n10 , \oc8051_top_1/oc8051_decoder1/n303 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n11 , \oc8051_top_1/oc8051_decoder1/n307 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n10 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n11 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n13 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n14 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n740 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n15 , \oc8051_top_1/oc8051_decoder1/n750 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n14 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n15 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_551/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n16 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n552 , \oc8051_top_1/oc8051_decoder1/reduce_or_551/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_551/n17 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_552/n2 , \oc8051_top_1/oc8051_decoder1/n217 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_552/n3 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_552/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n553 , \oc8051_top_1/oc8051_decoder1/reduce_or_552/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_552/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n2 , \oc8051_top_1/oc8051_decoder1/n543 , 
        \oc8051_top_1/oc8051_decoder1/n539 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n4 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n5 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/n86 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n6 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n5 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n7 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n9 , \oc8051_top_1/oc8051_decoder1/n512 , 
        \oc8051_top_1/oc8051_decoder1/n509 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n10 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/n497 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n11 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n10 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n11 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n13 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n490 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n14 , \oc8051_top_1/oc8051_decoder1/n482 , 
        \oc8051_top_1/oc8051_decoder1/n477 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n15 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n14 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n15 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n16 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n17 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n19 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n20 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n456 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n21 , \oc8051_top_1/oc8051_decoder1/n464 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n20 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n21 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n23 , \oc8051_top_1/oc8051_decoder1/n452 , 
        \oc8051_top_1/oc8051_decoder1/n446 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n24 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n25 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n24 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n25 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n26 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n28 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n936 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n29 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n922 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n30 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n29 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n30 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n32 , \oc8051_top_1/oc8051_decoder1/n402 , 
        \oc8051_top_1/oc8051_decoder1/n397 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n33 , \oc8051_top_1/oc8051_decoder1/n107 , 
        \oc8051_top_1/oc8051_decoder1/n382 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n34 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n33 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n34 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n35 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n37 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n36 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n38 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n37 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n39 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n861 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n40 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n41 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n39 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n40 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n42 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n839 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n43 , \oc8051_top_1/oc8051_decoder1/n348 , 
        \oc8051_top_1/oc8051_decoder1/n822 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n44 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n43 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n45 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n42 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n44 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n46 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n41 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n45 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n47 , \oc8051_top_1/oc8051_decoder1/n816 , 
        \oc8051_top_1/oc8051_decoder1/n811 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n48 , \oc8051_top_1/oc8051_decoder1/n323 , 
        \oc8051_top_1/oc8051_decoder1/n317 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n49 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n48 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n50 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n47 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n49 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n51 , \oc8051_top_1/oc8051_decoder1/n312 , 
        \oc8051_top_1/oc8051_decoder1/n307 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n52 , \oc8051_top_1/oc8051_decoder1/n763 , 
        \oc8051_top_1/oc8051_decoder1/n760 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n53 , \oc8051_top_1/oc8051_decoder1/n303 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n52 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n54 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n51 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n53 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n55 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n50 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n54 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n56 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n46 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n55 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n57 , \oc8051_top_1/oc8051_decoder1/n101 , 
        \oc8051_top_1/oc8051_decoder1/n750 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n58 , \oc8051_top_1/oc8051_decoder1/n740 , 
        \oc8051_top_1/oc8051_decoder1/n270 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n59 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n58 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n60 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n57 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n59 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n61 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n62 , \oc8051_top_1/oc8051_decoder1/n255 , 
        \oc8051_top_1/oc8051_decoder1/n252 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n63 , \oc8051_top_1/oc8051_decoder1/n258 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n62 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n64 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n61 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n63 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n65 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n60 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n64 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n66 , \oc8051_top_1/oc8051_decoder1/n248 , 
        \oc8051_top_1/oc8051_decoder1/n698 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n67 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n68 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n67 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n69 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n66 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n68 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n70 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/n679 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n71 , \oc8051_top_1/oc8051_decoder1/n217 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n72 , \oc8051_top_1/oc8051_decoder1/n675 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n71 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n73 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n70 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n72 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n74 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n69 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n73 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n75 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n65 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n74 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_554/n76 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n75 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n555 , \oc8051_top_1/oc8051_decoder1/reduce_or_554/n38 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_554/n76 ) ;   // oc8051_decoder.v(1223)
    and (\oc8051_top_1/oc8051_decoder1/Select_556/n2 , 1'b1, \oc8051_top_1/oc8051_decoder1/n556 ) ;   // oc8051_decoder.v(1223)
    and (\oc8051_top_1/oc8051_decoder1/Select_556/n3 , 1'b0, \oc8051_top_1/oc8051_decoder1/n555 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/Select_556/n4 , \oc8051_top_1/oc8051_decoder1/Select_556/n2 , 
        \oc8051_top_1/oc8051_decoder1/Select_556/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n557 , \oc8051_top_1/oc8051_decoder1/Select_556/n1 , 
        \oc8051_top_1/oc8051_decoder1/Select_556/n4 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_557/n2 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n425 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_557/n3 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_557/n2 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n558 , \oc8051_top_1/oc8051_decoder1/reduce_or_557/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_557/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n559 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_558/n1 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n2 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n1 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n3 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/n505 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n4 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/n497 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n4 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n5 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n7 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n490 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n8 , \oc8051_top_1/oc8051_decoder1/n936 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n8 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n10 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n402 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n11 , \oc8051_top_1/oc8051_decoder1/n397 , 
        \oc8051_top_1/oc8051_decoder1/n382 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n11 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n12 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n13 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n15 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n861 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n16 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n16 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n18 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n348 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n19 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n19 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n20 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n22 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n750 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n23 , \oc8051_top_1/oc8051_decoder1/n270 , 
        \oc8051_top_1/oc8051_decoder1/n258 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n23 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n25 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/n241 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n26 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n683 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n26 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n28 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n27 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_559/n29 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n28 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n560 , \oc8051_top_1/oc8051_decoder1/reduce_or_559/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_559/n29 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n2 , \oc8051_top_1/oc8051_decoder1/n199 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n1 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n3 , \oc8051_top_1/oc8051_decoder1/n477 , 
        \oc8051_top_1/oc8051_decoder1/n473 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n4 , \oc8051_top_1/oc8051_decoder1/n482 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n4 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n6 , \oc8051_top_1/oc8051_decoder1/n446 , 
        _cvpt_41) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n7 , \oc8051_top_1/oc8051_decoder1/n469 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n8 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/n433 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n9 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n8 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n9 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n10 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n12 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n13 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n12 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n14 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n15 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n14 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n15 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n17 , \oc8051_top_1/oc8051_decoder1/n317 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n18 , \oc8051_top_1/oc8051_decoder1/n323 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n17 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n19 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n20 , \oc8051_top_1/oc8051_decoder1/n217 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n20 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n21 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_560/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n22 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n561 , \oc8051_top_1/oc8051_decoder1/reduce_or_560/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_560/n23 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n2 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n1 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n3 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n436 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n4 , \oc8051_top_1/oc8051_decoder1/n464 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n3 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n4 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n6 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n402 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n7 , \oc8051_top_1/oc8051_decoder1/n127 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n6 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n8 , \oc8051_top_1/oc8051_decoder1/n382 , 
        \oc8051_top_1/oc8051_decoder1/n378 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n9 , \oc8051_top_1/oc8051_decoder1/n397 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n8 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_563/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n9 ) ;   // oc8051_decoder.v(1223)
    or (\oc8051_top_1/oc8051_decoder1/n564 , \oc8051_top_1/oc8051_decoder1/reduce_or_563/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_563/n10 ) ;   // oc8051_decoder.v(1223)
    assign \oc8051_top_1/oc8051_decoder1/Mux_565/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n145 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/ram_rd_sel [2] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_565/n2  : \oc8051_top_1/oc8051_decoder1/Mux_565/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_566/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n209  : \oc8051_top_1/oc8051_decoder1/n146 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/ram_rd_sel [1] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_566/n2  : \oc8051_top_1/oc8051_decoder1/Mux_566/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_567/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n209  : \oc8051_top_1/oc8051_decoder1/n147 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/ram_rd_sel [0] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_567/n2  : \oc8051_top_1/oc8051_decoder1/Mux_567/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_568/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n209  : \oc8051_top_1/oc8051_decoder1/n152 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/pc_wr  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_568/n2  : \oc8051_top_1/oc8051_decoder1/Mux_568/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_569/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n433 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/pc_wr_sel [2] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_569/n2  : \oc8051_top_1/oc8051_decoder1/Mux_569/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_570/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n154 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/pc_wr_sel [1] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_570/n2  : \oc8051_top_1/oc8051_decoder1/Mux_570/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_571/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n209  : \oc8051_top_1/oc8051_decoder1/n155 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/pc_wr_sel [0] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_571/n2  : \oc8051_top_1/oc8051_decoder1/Mux_571/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_572/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n199  : 1'b0;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/leave_su_mode  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_572/n2  : \oc8051_top_1/oc8051_decoder1/Mux_572/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_573/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n156 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/comp_sel [1] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_573/n2  : \oc8051_top_1/oc8051_decoder1/Mux_573/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_574/n2  = _cvpt_40 ? 1'b1 : \oc8051_top_1/oc8051_decoder1/n158 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/comp_sel [0] = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_574/n2  : \oc8051_top_1/oc8051_decoder1/Mux_574/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_575/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/rmw  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_575/n2  : \oc8051_top_1/oc8051_decoder1/Mux_575/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_576/n2  = _cvpt_40 ? 1'b1 : 1'b1;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/stb_i  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_576/n2  : \oc8051_top_1/oc8051_decoder1/Mux_576/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_577/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n159 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/bit_addr  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_577/n2  : \oc8051_top_1/oc8051_decoder1/Mux_577/n1 ;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/oc8051_decoder1/Mux_578/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(1225)
    assign \oc8051_top_1/enter_su_mode  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_578/n2  : \oc8051_top_1/oc8051_decoder1/Mux_578/n1 ;   // oc8051_decoder.v(1225)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_606/n2 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n1 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_606/n3 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_606/n4 , \oc8051_top_1/oc8051_decoder1/n477 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n3 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_606/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n4 ) ;   // oc8051_decoder.v(1347)
    not (\oc8051_top_1/oc8051_decoder1/n607 , \oc8051_top_1/oc8051_decoder1/reduce_nor_606/n5 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/n611 , \oc8051_top_1/oc8051_decoder1/n607 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_610/n1 ) ;   // oc8051_decoder.v(1347)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_639/n2 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n1 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_639/n3 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_639/n4 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n3 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_639/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n4 ) ;   // oc8051_decoder.v(1411)
    not (\oc8051_top_1/oc8051_decoder1/n640 , \oc8051_top_1/oc8051_decoder1/reduce_nor_639/n5 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/n641 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/reduce_or_640/n1 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/n642 , \oc8051_top_1/oc8051_decoder1/n640 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_641/n1 ) ;   // oc8051_decoder.v(1411)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_708/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1568)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_708/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n2 ) ;   // oc8051_decoder.v(1568)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_708/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n3 ) ;   // oc8051_decoder.v(1568)
    not (\oc8051_top_1/oc8051_decoder1/n709 , \oc8051_top_1/oc8051_decoder1/reduce_nor_708/n4 ) ;   // oc8051_decoder.v(1568)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_717/n2 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1590)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_717/n3 , \oc8051_top_1/oc8051_decoder1/n56 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n2 ) ;   // oc8051_decoder.v(1590)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_717/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n3 ) ;   // oc8051_decoder.v(1590)
    not (\oc8051_top_1/oc8051_decoder1/n718 , \oc8051_top_1/oc8051_decoder1/reduce_nor_717/n4 ) ;   // oc8051_decoder.v(1590)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n1 ) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n4 ) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_779/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n5 ) ;   // oc8051_decoder.v(1746)
    not (\oc8051_top_1/oc8051_decoder1/n780 , \oc8051_top_1/oc8051_decoder1/reduce_nor_779/n6 ) ;   // oc8051_decoder.v(1746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n2 , \oc8051_top_1/oc8051_decoder1/n84 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n1 ) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n3 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n4 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n4 ) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_790/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n5 ) ;   // oc8051_decoder.v(1768)
    not (\oc8051_top_1/oc8051_decoder1/n791 , \oc8051_top_1/oc8051_decoder1/reduce_nor_790/n6 ) ;   // oc8051_decoder.v(1768)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n2 ) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n5 ) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_833/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n6 ) ;   // oc8051_decoder.v(1869)
    not (\oc8051_top_1/oc8051_decoder1/n834 , \oc8051_top_1/oc8051_decoder1/reduce_nor_833/n7 ) ;   // oc8051_decoder.v(1869)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n2 ) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n5 ) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_842/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n6 ) ;   // oc8051_decoder.v(1891)
    not (\oc8051_top_1/oc8051_decoder1/n843 , \oc8051_top_1/oc8051_decoder1/reduce_nor_842/n7 ) ;   // oc8051_decoder.v(1891)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n2 ) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n5 ) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_883/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n6 ) ;   // oc8051_decoder.v(1990)
    not (\oc8051_top_1/oc8051_decoder1/n884 , \oc8051_top_1/oc8051_decoder1/reduce_nor_883/n7 ) ;   // oc8051_decoder.v(1990)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n2 ) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n5 ) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_888/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n6 ) ;   // oc8051_decoder.v(2001)
    not (\oc8051_top_1/oc8051_decoder1/n889 , \oc8051_top_1/oc8051_decoder1/reduce_nor_888/n7 ) ;   // oc8051_decoder.v(2001)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n2 ) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n5 ) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_898/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n6 ) ;   // oc8051_decoder.v(2023)
    not (\oc8051_top_1/oc8051_decoder1/n899 , \oc8051_top_1/oc8051_decoder1/reduce_nor_898/n7 ) ;   // oc8051_decoder.v(2023)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n2 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n5 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_904/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n6 ) ;   // oc8051_decoder.v(2034)
    not (\oc8051_top_1/oc8051_decoder1/n905 , \oc8051_top_1/oc8051_decoder1/reduce_nor_904/n7 ) ;   // oc8051_decoder.v(2034)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n2 ) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n5 ) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_914/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n6 ) ;   // oc8051_decoder.v(2056)
    not (\oc8051_top_1/oc8051_decoder1/n915 , \oc8051_top_1/oc8051_decoder1/reduce_nor_914/n7 ) ;   // oc8051_decoder.v(2056)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n2 ) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n5 ) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_917/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n6 ) ;   // oc8051_decoder.v(2067)
    not (\oc8051_top_1/oc8051_decoder1/n918 , \oc8051_top_1/oc8051_decoder1/reduce_nor_917/n7 ) ;   // oc8051_decoder.v(2067)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n2 ) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n5 ) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_932/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n6 ) ;   // oc8051_decoder.v(2111)
    not (\oc8051_top_1/oc8051_decoder1/n933 , \oc8051_top_1/oc8051_decoder1/reduce_nor_932/n7 ) ;   // oc8051_decoder.v(2111)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n2 ) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n5 ) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_986/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n6 ) ;   // oc8051_decoder.v(2278)
    not (\oc8051_top_1/oc8051_decoder1/n987 , \oc8051_top_1/oc8051_decoder1/reduce_nor_986/n7 ) ;   // oc8051_decoder.v(2278)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n2 ) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n5 ) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_993/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n6 ) ;   // oc8051_decoder.v(2289)
    not (\oc8051_top_1/oc8051_decoder1/n994 , \oc8051_top_1/oc8051_decoder1/reduce_nor_993/n7 ) ;   // oc8051_decoder.v(2289)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n2 ) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n5 ) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n6 ) ;   // oc8051_decoder.v(2311)
    not (\oc8051_top_1/oc8051_decoder1/n1004 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1003/n7 ) ;   // oc8051_decoder.v(2311)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n2 ) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n5 ) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n6 ) ;   // oc8051_decoder.v(2344)
    not (\oc8051_top_1/oc8051_decoder1/n1015 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1014/n7 ) ;   // oc8051_decoder.v(2344)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n2 ) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n5 ) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n6 ) ;   // oc8051_decoder.v(2421)
    not (\oc8051_top_1/oc8051_decoder1/n1044 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1043/n7 ) ;   // oc8051_decoder.v(2421)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n2 ) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n5 ) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n6 ) ;   // oc8051_decoder.v(2520)
    not (\oc8051_top_1/oc8051_decoder1/n1077 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1076/n7 ) ;   // oc8051_decoder.v(2520)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n2 ) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n5 ) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n6 ) ;   // oc8051_decoder.v(2531)
    not (\oc8051_top_1/oc8051_decoder1/n1082 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1081/n7 ) ;   // oc8051_decoder.v(2531)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n2 ) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n5 ) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n6 ) ;   // oc8051_decoder.v(2542)
    not (\oc8051_top_1/oc8051_decoder1/n1085 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1084/n7 ) ;   // oc8051_decoder.v(2542)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n2 ) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n5 ) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n6 ) ;   // oc8051_decoder.v(2553)
    not (\oc8051_top_1/oc8051_decoder1/n1089 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1088/n7 ) ;   // oc8051_decoder.v(2553)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n2 , \oc8051_top_1/op1_cur [2], 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n2 ) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n5 ) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n6 ) ;   // oc8051_decoder.v(2564)
    not (\oc8051_top_1/oc8051_decoder1/n1095 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1094/n7 ) ;   // oc8051_decoder.v(2564)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n2 ) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n4 , \oc8051_top_1/oc8051_decoder1/n74 , 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n5 , \oc8051_top_1/op1_d [6], 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n5 ) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n6 ) ;   // oc8051_decoder.v(2608)
    not (\oc8051_top_1/oc8051_decoder1/n1111 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1110/n7 ) ;   // oc8051_decoder.v(2608)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n2 ) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/op1_d [5]) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/oc8051_decoder1/n53 ) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n5 ) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n6 ) ;   // oc8051_decoder.v(2619)
    not (\oc8051_top_1/oc8051_decoder1/n1115 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1114/n7 ) ;   // oc8051_decoder.v(2619)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n2 , \oc8051_top_1/oc8051_decoder1/n52 , 
        \oc8051_top_1/op1_d [3]) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n2 ) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n4 , \oc8051_top_1/op1_d [4], 
        \oc8051_top_1/oc8051_decoder1/n56 ) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n5 , \oc8051_top_1/oc8051_decoder1/n72 , 
        \oc8051_top_1/op1_d [7]) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n5 ) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n6 ) ;   // oc8051_decoder.v(2652)
    not (\oc8051_top_1/oc8051_decoder1/n1129 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1128/n7 ) ;   // oc8051_decoder.v(2652)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n2 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n3 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n3 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n5 , \oc8051_top_1/oc8051_decoder1/n312 , 
        \oc8051_top_1/oc8051_decoder1/n780 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n6 , \oc8051_top_1/oc8051_decoder1/n791 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n7 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n8 , \oc8051_top_1/oc8051_decoder1/n763 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1139/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n8 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1140 , \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1139/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n2 , \oc8051_top_1/oc8051_decoder1/n548 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n3 , \oc8051_top_1/oc8051_decoder1/n512 , 
        \oc8051_top_1/oc8051_decoder1/n509 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n4 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n3 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n6 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n464 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n7 , \oc8051_top_1/oc8051_decoder1/n497 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n8 , \oc8051_top_1/oc8051_decoder1/n456 , 
        \oc8051_top_1/oc8051_decoder1/n994 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n9 , \oc8051_top_1/oc8051_decoder1/n1004 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n8 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n12 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/n936 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n13 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n14 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n402 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n15 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n17 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n18 , \oc8051_top_1/oc8051_decoder1/n397 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n19 , \oc8051_top_1/oc8051_decoder1/n255 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n20 , \oc8051_top_1/oc8051_decoder1/n307 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n19 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1140/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1141 , \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1140/n22 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1141/n2 , \oc8051_top_1/oc8051_decoder1/n439 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1142 , \oc8051_top_1/oc8051_decoder1/reduce_or_1141/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1141/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n2 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n4 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1085 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n5 , \oc8051_top_1/oc8051_decoder1/n1077 , 
        \oc8051_top_1/oc8051_decoder1/n497 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n6 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n9 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n10 , \oc8051_top_1/oc8051_decoder1/n1004 , 
        \oc8051_top_1/oc8051_decoder1/n994 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n11 , \oc8051_top_1/oc8051_decoder1/n1015 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n13 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n933 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n14 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/n915 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n15 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n16 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n19 , \oc8051_top_1/oc8051_decoder1/n899 , 
        \oc8051_top_1/oc8051_decoder1/n884 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n20 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n22 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n23 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n831 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n24 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n27 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n780 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n28 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n740 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n29 , \oc8051_top_1/oc8051_decoder1/n750 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n28 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n31 , \oc8051_top_1/oc8051_decoder1/n728 , 
        \oc8051_top_1/oc8051_decoder1/n709 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n32 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/n675 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n33 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n33 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n34 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1142/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n35 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1143 , \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1142/n36 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n2 , \oc8051_top_1/oc8051_decoder1/n1107 , 
        \oc8051_top_1/oc8051_decoder1/n1089 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n3 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n4 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n3 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n5 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/n1077 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n6 , \oc8051_top_1/oc8051_decoder1/n1085 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n7 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n473 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n8 , \oc8051_top_1/oc8051_decoder1/n1044 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n9 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n8 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n11 , \oc8051_top_1/oc8051_decoder1/n469 , 
        \oc8051_top_1/oc8051_decoder1/n994 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n12 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/n439 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n13 , \oc8051_top_1/oc8051_decoder1/n987 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n13 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n15 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n16 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n17 , \oc8051_top_1/oc8051_decoder1/n915 , 
        \oc8051_top_1/oc8051_decoder1/n899 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n18 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n18 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n20 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n19 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n22 , \oc8051_top_1/oc8051_decoder1/n884 , 
        \oc8051_top_1/oc8051_decoder1/n112 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n23 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n24 , \oc8051_top_1/oc8051_decoder1/n107 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n26 , \oc8051_top_1/oc8051_decoder1/n843 , 
        \oc8051_top_1/oc8051_decoder1/n839 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n27 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n26 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n28 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/n811 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n29 , \oc8051_top_1/oc8051_decoder1/n834 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n28 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n30 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n32 , \oc8051_top_1/oc8051_decoder1/n780 , 
        \oc8051_top_1/oc8051_decoder1/n750 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n33 , \oc8051_top_1/oc8051_decoder1/n791 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n34 , \oc8051_top_1/oc8051_decoder1/n740 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n35 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n34 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n33 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n35 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n37 , \oc8051_top_1/oc8051_decoder1/n709 , 
        \oc8051_top_1/oc8051_decoder1/n683 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n38 , \oc8051_top_1/oc8051_decoder1/n718 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n37 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n39 , \oc8051_top_1/oc8051_decoder1/n675 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n40 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n39 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n41 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n38 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n40 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n42 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n36 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n41 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1143/n43 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n42 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1144 , \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1143/n43 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n2 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n936 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n4 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n5 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n918 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n8 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n9 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n11 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/n241 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n12 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1144/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n13 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1145 , \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1144/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n2 , \oc8051_top_1/oc8051_decoder1/n543 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n3 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n493 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n4 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n3 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n6 , \oc8051_top_1/oc8051_decoder1/n490 , 
        \oc8051_top_1/oc8051_decoder1/n473 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n7 , \oc8051_top_1/oc8051_decoder1/n1044 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n8 , \oc8051_top_1/oc8051_decoder1/n884 , 
        \oc8051_top_1/oc8051_decoder1/n112 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n9 , \oc8051_top_1/oc8051_decoder1/n1015 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n8 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n12 , \oc8051_top_1/oc8051_decoder1/n843 , 
        \oc8051_top_1/oc8051_decoder1/n834 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n13 , \oc8051_top_1/oc8051_decoder1/n852 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n14 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n15 , \oc8051_top_1/oc8051_decoder1/n348 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n17 , \oc8051_top_1/oc8051_decoder1/n101 , 
        \oc8051_top_1/oc8051_decoder1/n270 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n18 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n19 , \oc8051_top_1/oc8051_decoder1/n258 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n20 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n19 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1145/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1146 , \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1145/n22 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n2 , \oc8051_top_1/oc8051_decoder1/n1129 , 
        \oc8051_top_1/oc8051_decoder1/n539 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n4 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n1115 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n5 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1085 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n8 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/n1077 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n9 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/n502 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n11 , \oc8051_top_1/oc8051_decoder1/n497 , 
        \oc8051_top_1/oc8051_decoder1/n493 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n12 , \oc8051_top_1/oc8051_decoder1/n490 , 
        \oc8051_top_1/oc8051_decoder1/n936 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n13 , \oc8051_top_1/oc8051_decoder1/n1044 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n13 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n17 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n18 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n918 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n18 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n20 , \oc8051_top_1/oc8051_decoder1/n382 , 
        \oc8051_top_1/oc8051_decoder1/n348 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n21 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n22 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n24 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n25 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n270 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n27 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n258 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n28 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/n691 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n29 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n28 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n30 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1146/n32 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n31 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1147 , \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1146/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n3 , \oc8051_top_1/oc8051_decoder1/n936 , 
        \oc8051_top_1/oc8051_decoder1/n933 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n4 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/n139 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n7 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/n915 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n8 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n9 , \oc8051_top_1/oc8051_decoder1/n402 , 
        \oc8051_top_1/oc8051_decoder1/n905 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n10 , \oc8051_top_1/oc8051_decoder1/n899 , 
        \oc8051_top_1/oc8051_decoder1/n382 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n14 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n15 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n16 , \oc8051_top_1/oc8051_decoder1/n852 , 
        \oc8051_top_1/oc8051_decoder1/n848 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n17 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n18 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n20 , \oc8051_top_1/oc8051_decoder1/n763 , 
        \oc8051_top_1/oc8051_decoder1/n760 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n21 , \oc8051_top_1/oc8051_decoder1/n750 , 
        \oc8051_top_1/oc8051_decoder1/n732 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n23 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/n241 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n24 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n683 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1147/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n26 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1148 , \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1147/n27 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n2 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n4 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/n1077 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n5 , \oc8051_top_1/oc8051_decoder1/n143 , 
        \oc8051_top_1/oc8051_decoder1/n936 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n6 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n9 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n10 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/n402 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n11 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n13 , \oc8051_top_1/oc8051_decoder1/n905 , 
        \oc8051_top_1/oc8051_decoder1/n899 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n14 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n15 , \oc8051_top_1/oc8051_decoder1/n884 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n16 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n19 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n861 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n20 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n22 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n822 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n23 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n24 , \oc8051_top_1/oc8051_decoder1/n816 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n27 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n101 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n28 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n29 , \oc8051_top_1/oc8051_decoder1/n750 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n28 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n31 , \oc8051_top_1/oc8051_decoder1/n698 , 
        \oc8051_top_1/oc8051_decoder1/n241 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n32 , \oc8051_top_1/oc8051_decoder1/n95 , 
        \oc8051_top_1/oc8051_decoder1/n683 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n33 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n33 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n34 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1148/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n35 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1149 , \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1148/n36 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n2 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1082 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n4 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/n497 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n5 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n1044 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n8 , \oc8051_top_1/oc8051_decoder1/n490 , 
        \oc8051_top_1/oc8051_decoder1/n143 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n9 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n469 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n11 , \oc8051_top_1/oc8051_decoder1/n433 , 
        \oc8051_top_1/oc8051_decoder1/n941 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n12 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n861 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n13 , \oc8051_top_1/oc8051_decoder1/n915 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n14 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n13 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n15 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n17 , \oc8051_top_1/oc8051_decoder1/n856 , 
        \oc8051_top_1/oc8051_decoder1/n852 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n18 , \oc8051_top_1/oc8051_decoder1/n848 , 
        \oc8051_top_1/oc8051_decoder1/n843 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n18 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n20 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n834 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n21 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n22 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n22 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n25 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/n750 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n26 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n740 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n25 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n26 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n28 , \oc8051_top_1/oc8051_decoder1/n732 , 
        \oc8051_top_1/oc8051_decoder1/n258 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n29 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/n675 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n30 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n30 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n32 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n31 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1149/n33 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1150 , \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1149/n33 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/n524 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n4 , \oc8051_top_1/oc8051_decoder1/n512 , 
        \oc8051_top_1/oc8051_decoder1/n509 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n5 , \oc8051_top_1/oc8051_decoder1/n493 , 
        \oc8051_top_1/oc8051_decoder1/n464 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n6 , \oc8051_top_1/oc8051_decoder1/n497 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n9 , \oc8051_top_1/oc8051_decoder1/n1004 , 
        \oc8051_top_1/oc8051_decoder1/n456 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n10 , _cvpt_41, \oc8051_top_1/oc8051_decoder1/n439 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n11 , \oc8051_top_1/oc8051_decoder1/n994 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n13 , \oc8051_top_1/oc8051_decoder1/n936 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n14 , \oc8051_top_1/oc8051_decoder1/n402 , 
        \oc8051_top_1/oc8051_decoder1/n397 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n15 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n16 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n19 , \oc8051_top_1/oc8051_decoder1/n861 , 
        \oc8051_top_1/oc8051_decoder1/n856 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n20 , \oc8051_top_1/oc8051_decoder1/n822 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n22 , \oc8051_top_1/oc8051_decoder1/n791 , 
        \oc8051_top_1/oc8051_decoder1/n312 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n23 , \oc8051_top_1/oc8051_decoder1/n307 , 
        \oc8051_top_1/oc8051_decoder1/n763 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n24 , \oc8051_top_1/oc8051_decoder1/n780 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n27 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n732 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n28 , \oc8051_top_1/oc8051_decoder1/n718 , 
        \oc8051_top_1/oc8051_decoder1/n252 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n29 , \oc8051_top_1/oc8051_decoder1/n255 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n28 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n30 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n31 , \oc8051_top_1/oc8051_decoder1/n709 , 
        \oc8051_top_1/oc8051_decoder1/n698 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n32 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n215 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n33 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n32 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n34 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n33 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n30 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n34 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1150/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n26 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n35 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1151 , \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1150/n36 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n2 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n3 , \oc8051_top_1/oc8051_decoder1/n139 , 
        \oc8051_top_1/oc8051_decoder1/n843 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n4 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n834 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n7 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n745 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n8 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n9 , \oc8051_top_1/oc8051_decoder1/n740 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n10 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/n675 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1151/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1152 , \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1151/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n2 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n3 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/n505 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n4 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n3 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n6 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n915 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n7 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n8 , \oc8051_top_1/oc8051_decoder1/n905 , 
        \oc8051_top_1/oc8051_decoder1/n889 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n9 , \oc8051_top_1/oc8051_decoder1/n112 , 
        \oc8051_top_1/oc8051_decoder1/n107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n9 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n13 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n843 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n14 , \oc8051_top_1/oc8051_decoder1/n382 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n13 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n15 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n834 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n16 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/n811 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n16 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n19 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n740 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n20 , \oc8051_top_1/oc8051_decoder1/n101 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n19 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n21 , \oc8051_top_1/oc8051_decoder1/n728 , 
        \oc8051_top_1/oc8051_decoder1/n95 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n22 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/n675 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n23 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n22 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n24 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n23 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1152/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1153 , \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1152/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n3 , \oc8051_top_1/oc8051_decoder1/n460 , 
        \oc8051_top_1/oc8051_decoder1/n941 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n4 , \oc8051_top_1/oc8051_decoder1/n415 , 
        \oc8051_top_1/oc8051_decoder1/n922 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n7 , \oc8051_top_1/oc8051_decoder1/n402 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n8 , \oc8051_top_1/oc8051_decoder1/n918 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n9 , \oc8051_top_1/oc8051_decoder1/n760 , 
        \oc8051_top_1/oc8051_decoder1/n732 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n10 , \oc8051_top_1/oc8051_decoder1/n241 , 
        \oc8051_top_1/oc8051_decoder1/n691 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1153/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1154 , \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1153/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n3 , \oc8051_top_1/oc8051_decoder1/n524 , 
        \oc8051_top_1/oc8051_decoder1/n1095 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n4 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1082 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n7 , \oc8051_top_1/oc8051_decoder1/n502 , 
        \oc8051_top_1/oc8051_decoder1/n464 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n8 , \oc8051_top_1/oc8051_decoder1/n505 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n9 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n415 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n10 , \oc8051_top_1/oc8051_decoder1/n922 , 
        \oc8051_top_1/oc8051_decoder1/n918 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n13 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n14 , \oc8051_top_1/oc8051_decoder1/n905 , 
        \oc8051_top_1/oc8051_decoder1/n382 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n15 , \oc8051_top_1/oc8051_decoder1/n915 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n16 , \oc8051_top_1/oc8051_decoder1/n378 , 
        \oc8051_top_1/oc8051_decoder1/n843 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n17 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n816 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n19 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n15 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n18 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n20 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/n760 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n21 , \oc8051_top_1/oc8051_decoder1/n745 , 
        \oc8051_top_1/oc8051_decoder1/n732 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n23 , \oc8051_top_1/oc8051_decoder1/n728 , 
        \oc8051_top_1/oc8051_decoder1/n241 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n24 , \oc8051_top_1/oc8051_decoder1/n691 , 
        \oc8051_top_1/oc8051_decoder1/n679 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n25 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1154/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n26 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1155 , \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1154/n27 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n2 , \oc8051_top_1/oc8051_decoder1/n71 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n3 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/n83 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n4 , \oc8051_top_1/oc8051_decoder1/n80 , 
        \oc8051_top_1/oc8051_decoder1/n76 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n6 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n7 , \oc8051_top_1/oc8051_decoder1/n73 , 
        \oc8051_top_1/oc8051_decoder1/n127 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n8 , \oc8051_top_1/oc8051_decoder1/n436 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n9 , \oc8051_top_1/oc8051_decoder1/n425 , 
        \oc8051_top_1/oc8051_decoder1/n397 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n10 , \oc8051_top_1/oc8051_decoder1/n889 , 
        \oc8051_top_1/oc8051_decoder1/n884 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1155/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1156 , \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1155/n12 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1156/n2 , \oc8051_top_1/oc8051_decoder1/n1120 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n1 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1156/n3 , \oc8051_top_1/oc8051_decoder1/n941 , 
        \oc8051_top_1/oc8051_decoder1/n822 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1156/n4 , \oc8051_top_1/oc8051_decoder1/n816 , 
        \oc8051_top_1/oc8051_decoder1/n732 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1156/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n4 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1157 , \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1156/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n2 , \oc8051_top_1/oc8051_decoder1/n1111 , 
        \oc8051_top_1/oc8051_decoder1/n1107 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n3 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n2 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n4 , \oc8051_top_1/oc8051_decoder1/n1089 , 
        \oc8051_top_1/oc8051_decoder1/n1085 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n5 , \oc8051_top_1/oc8051_decoder1/n1077 , 
        \oc8051_top_1/oc8051_decoder1/n1044 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n6 , \oc8051_top_1/oc8051_decoder1/n1082 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n5 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n7 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n6 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n8 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n7 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n9 , \oc8051_top_1/oc8051_decoder1/n490 , 
        \oc8051_top_1/oc8051_decoder1/n1015 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n10 , \oc8051_top_1/oc8051_decoder1/n452 , 
        \oc8051_top_1/oc8051_decoder1/n941 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n11 , \oc8051_top_1/oc8051_decoder1/n987 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n10 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n12 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n11 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n13 , \oc8051_top_1/oc8051_decoder1/n933 , 
        \oc8051_top_1/oc8051_decoder1/n918 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n14 , \oc8051_top_1/oc8051_decoder1/n899 , 
        \oc8051_top_1/oc8051_decoder1/n884 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n15 , \oc8051_top_1/oc8051_decoder1/n915 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n14 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n15 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n17 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n12 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n16 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n18 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n8 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n17 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n19 , \oc8051_top_1/oc8051_decoder1/n852 , 
        \oc8051_top_1/oc8051_decoder1/n848 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n20 , \oc8051_top_1/oc8051_decoder1/n839 , 
        \oc8051_top_1/oc8051_decoder1/n834 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n21 , \oc8051_top_1/oc8051_decoder1/n843 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n20 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n19 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n21 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n23 , \oc8051_top_1/oc8051_decoder1/n831 , 
        \oc8051_top_1/oc8051_decoder1/n348 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n24 , \oc8051_top_1/oc8051_decoder1/n327 , 
        \oc8051_top_1/oc8051_decoder1/n303 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n25 , \oc8051_top_1/oc8051_decoder1/n811 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n24 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n26 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n25 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n27 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n22 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n26 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n28 , \oc8051_top_1/oc8051_decoder1/n750 , 
        \oc8051_top_1/oc8051_decoder1/n745 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n29 , \oc8051_top_1/oc8051_decoder1/n270 , 
        \oc8051_top_1/oc8051_decoder1/n728 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n30 , \oc8051_top_1/oc8051_decoder1/n740 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n29 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n31 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n28 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n30 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n32 , \oc8051_top_1/oc8051_decoder1/n258 , 
        \oc8051_top_1/oc8051_decoder1/n248 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n33 , \oc8051_top_1/oc8051_decoder1/n679 , 
        \oc8051_top_1/oc8051_decoder1/n675 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n34 , \oc8051_top_1/oc8051_decoder1/n683 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n33 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n35 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n32 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n34 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n36 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n31 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n35 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1157/n37 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n27 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n36 ) ;   // oc8051_decoder.v(2696)
    or (\oc8051_top_1/oc8051_decoder1/n1158 , \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1157/n37 ) ;   // oc8051_decoder.v(2696)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1158/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n641 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1159  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1158/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1158/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1159/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n208 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1160  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1159/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1159/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1160/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n208 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1161  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1160/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1160/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1161/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1162  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1161/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1161/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1162/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1163  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1162/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1162/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1163/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1164  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1163/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1163/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1164/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n139  : \oc8051_top_1/oc8051_decoder1/n139 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1165  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1164/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1164/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1165/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n143  : \oc8051_top_1/oc8051_decoder1/n143 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1166  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1165/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1165/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1166/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n143  : \oc8051_top_1/oc8051_decoder1/n143 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1167  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1166/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1166/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1167/n2  = _cvpt_40 ? \oc8051_top_1/oc8051_decoder1/n208  : \oc8051_top_1/oc8051_decoder1/n208 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1168  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1167/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1167/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1168/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1169  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1168/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1168/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1169/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1170  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1169/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1169/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1170/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n641 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1171  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1170/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1170/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1171/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n643 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1172  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1171/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1171/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1172/n2  = _cvpt_40 ? 1'b0 : \oc8051_top_1/oc8051_decoder1/n643 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1173  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1172/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1172/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1173/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1174  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1173/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1173/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1174/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1175  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1174/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1174/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1175/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1176  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1175/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1175/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1176/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1177  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1176/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1176/n1 ;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1177/n2  = _cvpt_40 ? 1'b0 : 1'b0;   // oc8051_decoder.v(2698)
    assign \oc8051_top_1/oc8051_decoder1/n1178  = _cvpt_208 ? \oc8051_top_1/oc8051_decoder1/Mux_1177/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1177/n1 ;   // oc8051_decoder.v(2698)
    not (_cvpt_95, \oc8051_top_1/oc8051_decoder1/reduce_nor_1219/n1 ) ;   // oc8051_decoder.v(2707)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n2 , \oc8051_top_1/op1_n [3], 
        \oc8051_top_1/oc8051_decoder1/n1242 ) ;   // oc8051_decoder.v(2721)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n3 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n2 ) ;   // oc8051_decoder.v(2721)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n3 ) ;   // oc8051_decoder.v(2721)
    not (\oc8051_top_1/oc8051_decoder1/n1243 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1242/n4 ) ;   // oc8051_decoder.v(2721)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n2 , \oc8051_top_1/op1_n [3], 
        \oc8051_top_1/op1_n [4]) ;   // oc8051_decoder.v(2722)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n3 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n2 ) ;   // oc8051_decoder.v(2722)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n3 ) ;   // oc8051_decoder.v(2722)
    not (\oc8051_top_1/oc8051_decoder1/n1245 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1244/n4 ) ;   // oc8051_decoder.v(2722)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n2 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n3 , \oc8051_top_1/oc8051_decoder1/n1248 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n2 ) ;   // oc8051_decoder.v(2723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n3 ) ;   // oc8051_decoder.v(2723)
    not (\oc8051_top_1/oc8051_decoder1/n1250 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1249/n4 ) ;   // oc8051_decoder.v(2723)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n2 , \oc8051_top_1/oc8051_decoder1/n1251 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n1 ) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n3 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n4 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n4 ) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n5 ) ;   // oc8051_decoder.v(2724)
    not (\oc8051_top_1/oc8051_decoder1/n1256 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1255/n6 ) ;   // oc8051_decoder.v(2724)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n2 ) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n5 ) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n6 ) ;   // oc8051_decoder.v(2725)
    not (\oc8051_top_1/oc8051_decoder1/n1262 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1261/n7 ) ;   // oc8051_decoder.v(2725)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n2 ) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n5 ) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n6 ) ;   // oc8051_decoder.v(2726)
    not (\oc8051_top_1/oc8051_decoder1/n1267 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1266/n7 ) ;   // oc8051_decoder.v(2726)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n2 ) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n5 ) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n6 ) ;   // oc8051_decoder.v(2727)
    not (\oc8051_top_1/oc8051_decoder1/n1269 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1268/n7 ) ;   // oc8051_decoder.v(2727)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n2 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2728)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n3 , \oc8051_top_1/op1_n [5], 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n2 ) ;   // oc8051_decoder.v(2728)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n4 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n3 ) ;   // oc8051_decoder.v(2728)
    not (\oc8051_top_1/oc8051_decoder1/n1274 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1273/n4 ) ;   // oc8051_decoder.v(2728)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n2 ) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n5 ) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n6 ) ;   // oc8051_decoder.v(2729)
    not (\oc8051_top_1/oc8051_decoder1/n1280 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1279/n7 ) ;   // oc8051_decoder.v(2729)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n2 ) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n5 ) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n6 ) ;   // oc8051_decoder.v(2730)
    not (\oc8051_top_1/oc8051_decoder1/n1283 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1282/n7 ) ;   // oc8051_decoder.v(2730)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n2 ) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n5 ) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n6 ) ;   // oc8051_decoder.v(2731)
    not (\oc8051_top_1/oc8051_decoder1/n1288 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1287/n7 ) ;   // oc8051_decoder.v(2731)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n2 ) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n5 ) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n6 ) ;   // oc8051_decoder.v(2732)
    not (\oc8051_top_1/oc8051_decoder1/n1293 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1292/n7 ) ;   // oc8051_decoder.v(2732)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n2 ) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n5 ) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n6 ) ;   // oc8051_decoder.v(2733)
    not (\oc8051_top_1/oc8051_decoder1/n1297 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1296/n7 ) ;   // oc8051_decoder.v(2733)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n2 , \oc8051_top_1/oc8051_decoder1/n1251 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n1 ) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n3 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n4 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n4 ) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n5 ) ;   // oc8051_decoder.v(2734)
    not (\oc8051_top_1/oc8051_decoder1/n1302 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1301/n6 ) ;   // oc8051_decoder.v(2734)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n2 , \oc8051_top_1/oc8051_decoder1/n1251 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n1 ) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n3 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n4 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n4 ) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n5 ) ;   // oc8051_decoder.v(2735)
    not (\oc8051_top_1/oc8051_decoder1/n1308 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1307/n6 ) ;   // oc8051_decoder.v(2735)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n2 ) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n5 ) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n6 ) ;   // oc8051_decoder.v(2736)
    not (\oc8051_top_1/oc8051_decoder1/n1312 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1311/n7 ) ;   // oc8051_decoder.v(2736)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n2 ) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n5 ) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n6 ) ;   // oc8051_decoder.v(2737)
    not (\oc8051_top_1/oc8051_decoder1/n1317 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1316/n7 ) ;   // oc8051_decoder.v(2737)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n2 ) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n5 ) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n6 ) ;   // oc8051_decoder.v(2738)
    not (\oc8051_top_1/oc8051_decoder1/n1320 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1319/n7 ) ;   // oc8051_decoder.v(2738)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n2 ) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n5 ) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n6 ) ;   // oc8051_decoder.v(2739)
    not (\oc8051_top_1/oc8051_decoder1/n1324 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1323/n7 ) ;   // oc8051_decoder.v(2739)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n2 ) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n5 ) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n6 ) ;   // oc8051_decoder.v(2740)
    not (\oc8051_top_1/oc8051_decoder1/n1326 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1325/n7 ) ;   // oc8051_decoder.v(2740)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n2 ) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n5 ) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n6 ) ;   // oc8051_decoder.v(2741)
    not (\oc8051_top_1/oc8051_decoder1/n1328 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1327/n7 ) ;   // oc8051_decoder.v(2741)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n2 ) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n5 ) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n6 ) ;   // oc8051_decoder.v(2742)
    not (\oc8051_top_1/oc8051_decoder1/n1330 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1329/n7 ) ;   // oc8051_decoder.v(2742)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n2 ) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n5 ) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n6 ) ;   // oc8051_decoder.v(2743)
    not (\oc8051_top_1/oc8051_decoder1/n1332 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1331/n7 ) ;   // oc8051_decoder.v(2743)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n2 ) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n5 ) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n6 ) ;   // oc8051_decoder.v(2744)
    not (\oc8051_top_1/oc8051_decoder1/n1338 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1337/n7 ) ;   // oc8051_decoder.v(2744)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n2 ) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n5 ) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n6 ) ;   // oc8051_decoder.v(2745)
    not (\oc8051_top_1/oc8051_decoder1/n1341 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1340/n7 ) ;   // oc8051_decoder.v(2745)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n2 ) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n5 ) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n6 ) ;   // oc8051_decoder.v(2746)
    not (\oc8051_top_1/oc8051_decoder1/n1344 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1343/n7 ) ;   // oc8051_decoder.v(2746)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n2 ) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n4 , \oc8051_top_1/oc8051_decoder1/n1242 , 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n5 ) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n6 ) ;   // oc8051_decoder.v(2747)
    not (\oc8051_top_1/oc8051_decoder1/n1348 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1347/n7 ) ;   // oc8051_decoder.v(2747)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n2 , \oc8051_top_1/op1_n [2], 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n2 ) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n5 , \oc8051_top_1/oc8051_decoder1/n1272 , 
        \oc8051_top_1/op1_n [7]) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n5 ) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n6 ) ;   // oc8051_decoder.v(2748)
    not (\oc8051_top_1/oc8051_decoder1/n1351 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1350/n7 ) ;   // oc8051_decoder.v(2748)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n2 ) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/op1_n [5]) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n5 ) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n6 ) ;   // oc8051_decoder.v(2749)
    not (\oc8051_top_1/oc8051_decoder1/n1354 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1353/n7 ) ;   // oc8051_decoder.v(2749)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n2 , \oc8051_top_1/oc8051_decoder1/n1252 , 
        \oc8051_top_1/op1_n [3]) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n3 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n1 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n2 ) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n4 , \oc8051_top_1/op1_n [4], 
        \oc8051_top_1/oc8051_decoder1/n1248 ) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n5 , \oc8051_top_1/op1_n [6], 
        \oc8051_top_1/oc8051_decoder1/n1249 ) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n4 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n5 ) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n7 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n6 ) ;   // oc8051_decoder.v(2750)
    not (\oc8051_top_1/oc8051_decoder1/n1358 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1357/n7 ) ;   // oc8051_decoder.v(2750)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n2 , \oc8051_top_1/oc8051_decoder1/n1358 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n1 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n3 , \oc8051_top_1/oc8051_decoder1/n1348 , 
        \oc8051_top_1/oc8051_decoder1/n1344 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n4 , \oc8051_top_1/oc8051_decoder1/n1341 , 
        \oc8051_top_1/oc8051_decoder1/n1338 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n3 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n4 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n6 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n5 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n7 , \oc8051_top_1/oc8051_decoder1/n1332 , 
        \oc8051_top_1/oc8051_decoder1/n1330 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n8 , \oc8051_top_1/oc8051_decoder1/n1328 , 
        \oc8051_top_1/oc8051_decoder1/n1326 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n9 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n8 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n10 , \oc8051_top_1/oc8051_decoder1/n1324 , 
        \oc8051_top_1/oc8051_decoder1/n1320 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n11 , \oc8051_top_1/oc8051_decoder1/n1317 , 
        \oc8051_top_1/oc8051_decoder1/n1312 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n12 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n10 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n11 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n13 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n9 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n12 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n14 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n6 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n13 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n15 , \oc8051_top_1/oc8051_decoder1/n1302 , 
        \oc8051_top_1/oc8051_decoder1/n1297 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n16 , \oc8051_top_1/oc8051_decoder1/n1308 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n15 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n17 , \oc8051_top_1/oc8051_decoder1/n1293 , 
        \oc8051_top_1/oc8051_decoder1/n1288 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n18 , \oc8051_top_1/oc8051_decoder1/n1283 , 
        \oc8051_top_1/oc8051_decoder1/n1280 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n19 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n17 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n18 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n20 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n19 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n21 , \oc8051_top_1/oc8051_decoder1/n1274 , 
        \oc8051_top_1/oc8051_decoder1/n1269 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n22 , \oc8051_top_1/oc8051_decoder1/n1267 , 
        \oc8051_top_1/oc8051_decoder1/n1262 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n23 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n21 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n22 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n24 , \oc8051_top_1/oc8051_decoder1/n1256 , 
        \oc8051_top_1/oc8051_decoder1/n1250 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n25 , \oc8051_top_1/oc8051_decoder1/n1245 , 
        \oc8051_top_1/oc8051_decoder1/n1243 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n26 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n24 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n25 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n27 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n23 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n26 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n28 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n20 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n27 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n29 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n14 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n28 ) ;   // oc8051_decoder.v(2752)
    not (_cvpt_103, \oc8051_top_1/oc8051_decoder1/reduce_nor_1358/n29 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n2 , \oc8051_top_1/oc8051_decoder1/n1351 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n1 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n3 , \oc8051_top_1/oc8051_decoder1/n1338 , 
        \oc8051_top_1/oc8051_decoder1/n1332 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n4 , \oc8051_top_1/oc8051_decoder1/n1341 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n3 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n5 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n4 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n6 , \oc8051_top_1/oc8051_decoder1/n1328 , 
        \oc8051_top_1/oc8051_decoder1/n1326 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n7 , \oc8051_top_1/oc8051_decoder1/n1330 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n6 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n8 , \oc8051_top_1/oc8051_decoder1/n1312 , 
        \oc8051_top_1/oc8051_decoder1/n1308 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n9 , \oc8051_top_1/oc8051_decoder1/n1317 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n8 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n10 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n7 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n9 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n11 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n5 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n10 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n12 , \oc8051_top_1/oc8051_decoder1/n1288 , 
        \oc8051_top_1/oc8051_decoder1/n1283 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n13 , \oc8051_top_1/oc8051_decoder1/n1302 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n12 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n14 , \oc8051_top_1/oc8051_decoder1/n1274 , 
        \oc8051_top_1/oc8051_decoder1/n1269 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n15 , \oc8051_top_1/oc8051_decoder1/n1280 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n14 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n16 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n13 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n15 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n17 , \oc8051_top_1/oc8051_decoder1/n1262 , 
        \oc8051_top_1/oc8051_decoder1/n1256 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n18 , \oc8051_top_1/oc8051_decoder1/n1267 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n17 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n19 , \oc8051_top_1/oc8051_decoder1/n1245 , 
        \oc8051_top_1/oc8051_decoder1/n1243 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n20 , \oc8051_top_1/oc8051_decoder1/n1250 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n19 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n21 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n18 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n20 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1360/n22 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n16 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n21 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/n1361 , \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n11 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1360/n22 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1361/n2 , \oc8051_top_1/oc8051_decoder1/n1358 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n1 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1361/n3 , \oc8051_top_1/oc8051_decoder1/n1297 , 
        \oc8051_top_1/oc8051_decoder1/n1293 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/reduce_or_1361/n4 , \oc8051_top_1/oc8051_decoder1/n1320 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n3 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/n1362 , \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1361/n4 ) ;   // oc8051_decoder.v(2752)
    and (\oc8051_top_1/oc8051_decoder1/Select_1362/n2 , 1'b1, \oc8051_top_1/oc8051_decoder1/n1362 ) ;   // oc8051_decoder.v(2752)
    and (\oc8051_top_1/oc8051_decoder1/Select_1362/n3 , 1'b0, \oc8051_top_1/oc8051_decoder1/n1361 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/Select_1362/n4 , \oc8051_top_1/oc8051_decoder1/Select_1362/n2 , 
        \oc8051_top_1/oc8051_decoder1/Select_1362/n3 ) ;   // oc8051_decoder.v(2752)
    or (\oc8051_top_1/oc8051_decoder1/n1363 , \oc8051_top_1/oc8051_decoder1/Select_1362/n1 , 
        \oc8051_top_1/oc8051_decoder1/Select_1362/n4 ) ;   // oc8051_decoder.v(2752)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1363/n2  = _cvpt_104 ? 1'b1 : 1'b0;   // oc8051_decoder.v(2754)
    assign \oc8051_top_1/oc8051_decoder1/n1364  = _cvpt_276 ? \oc8051_top_1/oc8051_decoder1/Mux_1363/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1363/n1 ;   // oc8051_decoder.v(2754)
    assign \oc8051_top_1/oc8051_decoder1/Mux_1364/n2  = _cvpt_104 ? 1'b0 : 1'b1;   // oc8051_decoder.v(2754)
    assign \oc8051_top_1/oc8051_decoder1/n1365  = _cvpt_276 ? \oc8051_top_1/oc8051_decoder1/Mux_1364/n2  : \oc8051_top_1/oc8051_decoder1/Mux_1364/n1 ;   // oc8051_decoder.v(2754)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n2 , \oc8051_top_1/oc8051_decoder1/n473 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n1 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n3 , \oc8051_top_1/oc8051_decoder1/n482 , 
        \oc8051_top_1/oc8051_decoder1/n323 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n4 , \oc8051_top_1/oc8051_decoder1/n317 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n3 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n5 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n2 , 
        \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n4 ) ;   // oc8051_decoder.v(2785)
    not (\oc8051_top_1/oc8051_decoder1/n1418 , \oc8051_top_1/oc8051_decoder1/reduce_nor_1417/n5 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/n1419 , \oc8051_top_1/oc8051_decoder1/n1418 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1418/n1 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/n1420 , \oc8051_top_1/oc8051_decoder1/n1418 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1419/n1 ) ;   // oc8051_decoder.v(2785)
    or (\oc8051_top_1/oc8051_decoder1/n1421 , \oc8051_top_1/oc8051_decoder1/n1418 , 
        \oc8051_top_1/oc8051_decoder1/reduce_or_1420/n1 ) ;   // oc8051_decoder.v(2785)
    xor (_cvpt_3369, \oc8051_xiommu1/proc_addr [0], 1'b0) ;   // aes_top.v(94)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n1 , \oc8051_xiommu1/proc_addr [0], 
        \oc8051_xiommu1/proc_addr [1]) ;   // aes_top.v(97)
    and (\oc8051_xiommu1/aes_addr_range , \oc8051_xiommu1/aes_top_i/n4 , 
        \oc8051_xiommu1/aes_top_i/n5 ) ;   // aes_top.v(94)
    and (\oc8051_xiommu1/ack_aes , _cvpt_151, \oc8051_xiommu1/aes_addr_range ) ;   // aes_top.v(95)
    not (\oc8051_xiommu1/aes_top_i/n8 , \oc8051_xiommu1/proc_addr [8]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n9 , \oc8051_xiommu1/proc_addr [9]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n10 , \oc8051_xiommu1/proc_addr [10]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n11 , \oc8051_xiommu1/proc_addr [11]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n12 , \oc8051_xiommu1/proc_addr [12]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n13 , \oc8051_xiommu1/proc_addr [13]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n14 , \oc8051_xiommu1/proc_addr [14]) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/n15 , \oc8051_xiommu1/proc_addr [15]) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n1 , \oc8051_xiommu1/aes_top_i/n17 , 
        \oc8051_xiommu1/proc_addr [1]) ;   // aes_top.v(98)
    not (\oc8051_xiommu1/aes_top_i/n17 , \oc8051_xiommu1/proc_addr [0]) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n1 , \oc8051_xiommu1/proc_addr [0], 
        \oc8051_xiommu1/aes_top_i/n27 ) ;   // aes_top.v(99)
    not (\oc8051_xiommu1/aes_top_i/n27 , \oc8051_xiommu1/proc_addr [1]) ;   // aes_top.v(99)
    not (\oc8051_xiommu1/aes_top_i/n28 , \oc8051_xiommu1/proc_addr [2]) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n1 , \oc8051_xiommu1/proc_addr [2], 
        \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n1 , \oc8051_xiommu1/aes_top_i/n28 , 
        \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n1 , \oc8051_xiommu1/proc_addr [5], 
        \oc8051_xiommu1/proc_addr [6]) ;   // aes_top.v(102)
    not (\oc8051_xiommu1/aes_top_i/n58 , \oc8051_xiommu1/proc_addr [4]) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n1 , \oc8051_xiommu1/aes_top_i/n68 , 
        \oc8051_xiommu1/proc_addr [6]) ;   // aes_top.v(103)
    not (\oc8051_xiommu1/aes_top_i/n68 , \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n1 , \oc8051_xiommu1/aes_top_i/n68 , 
        \oc8051_xiommu1/proc_addr [6]) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_144/n1 , \oc8051_xiommu1/aes_state [0], 
        \oc8051_xiommu1/aes_state [1]) ;   // aes_top.v(120)
    assign \oc8051_xiommu1/aes_top_i/n89  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [7] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n90  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [6] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n91  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [5] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n92  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [4] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n93  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [3] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n94  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [2] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n95  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [1] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n96  = _cvpt_279 ? \oc8051_xiommu1/aes_top_i/aes_key1_dataout [0] : 1'b0;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n97  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [7] : \oc8051_xiommu1/aes_top_i/n89 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n98  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [6] : \oc8051_xiommu1/aes_top_i/n90 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n99  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [5] : \oc8051_xiommu1/aes_top_i/n91 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n100  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [4] : \oc8051_xiommu1/aes_top_i/n92 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n101  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [3] : \oc8051_xiommu1/aes_top_i/n93 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n102  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [2] : \oc8051_xiommu1/aes_top_i/n94 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n103  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [1] : \oc8051_xiommu1/aes_top_i/n95 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n104  = _cvpt_287 ? \oc8051_xiommu1/aes_top_i/aes_key0_dataout [0] : \oc8051_xiommu1/aes_top_i/n96 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n105  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [7] : \oc8051_xiommu1/aes_top_i/n97 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n106  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [6] : \oc8051_xiommu1/aes_top_i/n98 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n107  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [5] : \oc8051_xiommu1/aes_top_i/n99 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n108  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [4] : \oc8051_xiommu1/aes_top_i/n100 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n109  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [3] : \oc8051_xiommu1/aes_top_i/n101 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n110  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [2] : \oc8051_xiommu1/aes_top_i/n102 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n111  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [1] : \oc8051_xiommu1/aes_top_i/n103 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n112  = _cvpt_295 ? \oc8051_xiommu1/aes_top_i/aes_ctr_dataout [0] : \oc8051_xiommu1/aes_top_i/n104 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n113  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n105 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n114  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n106 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n115  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n107 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n116  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n108 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n117  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n109 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n118  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n110 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n119  = _cvpt_303 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n111 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n120  = _cvpt_303 ? _cvpt_538 : \oc8051_xiommu1/aes_top_i/n112 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n121  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [7] : \oc8051_xiommu1/aes_top_i/n113 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n122  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [6] : \oc8051_xiommu1/aes_top_i/n114 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n123  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [5] : \oc8051_xiommu1/aes_top_i/n115 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n124  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [4] : \oc8051_xiommu1/aes_top_i/n116 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n125  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [3] : \oc8051_xiommu1/aes_top_i/n117 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n126  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [2] : \oc8051_xiommu1/aes_top_i/n118 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n127  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [1] : \oc8051_xiommu1/aes_top_i/n119 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n128  = _cvpt_311 ? \oc8051_xiommu1/aes_top_i/aes_len_dataout [0] : \oc8051_xiommu1/aes_top_i/n120 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n129  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [7] : \oc8051_xiommu1/aes_top_i/n121 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n130  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [6] : \oc8051_xiommu1/aes_top_i/n122 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n131  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [5] : \oc8051_xiommu1/aes_top_i/n123 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n132  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [4] : \oc8051_xiommu1/aes_top_i/n124 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n133  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [3] : \oc8051_xiommu1/aes_top_i/n125 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n134  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [2] : \oc8051_xiommu1/aes_top_i/n126 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n135  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [1] : \oc8051_xiommu1/aes_top_i/n127 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/aes_top_i/n136  = _cvpt_319 ? \oc8051_xiommu1/aes_top_i/aes_addr_dataout [0] : \oc8051_xiommu1/aes_top_i/n128 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [7] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n129 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [6] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n130 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [5] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n131 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [4] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n132 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [3] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n133 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [2] = _cvpt_327 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n134 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [1] = _cvpt_327 ? \oc8051_xiommu1/aes_state [1] : \oc8051_xiommu1/aes_top_i/n135 ;   // aes_top.v(117)
    assign \oc8051_xiommu1/data_out_aes [0] = _cvpt_327 ? \oc8051_xiommu1/aes_state [0] : \oc8051_xiommu1/aes_top_i/n136 ;   // aes_top.v(117)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_146/n1 , \oc8051_xiommu1/aes_top_i/n146 , 
        \oc8051_xiommu1/aes_state [1]) ;   // aes_top.v(121)
    not (\oc8051_xiommu1/aes_top_i/n146 , \oc8051_xiommu1/aes_state [0]) ;   // aes_top.v(121)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_148/n1 , \oc8051_xiommu1/aes_state [0], 
        \oc8051_xiommu1/aes_top_i/n148 ) ;   // aes_top.v(122)
    not (\oc8051_xiommu1/aes_top_i/n148 , \oc8051_xiommu1/aes_state [1]) ;   // aes_top.v(122)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_151/n1 , \oc8051_xiommu1/aes_top_i/n146 , 
        \oc8051_xiommu1/aes_top_i/n148 ) ;   // aes_top.v(123)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [4]), 
            .b(1'b1), .o(\oc8051_xiommu1/aes_top_i/n176 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n2 ));   // aes_top.v(214)
    and (\oc8051_xiommu1/aes_top_i/wren , \oc8051_xiommu1/write_aes , _cvpt_408) ;   // aes_top.v(126)
    and (\oc8051_xiommu1/aes_top_i/n154 , \oc8051_xiommu1/aes_top_i/sel_reg_start , 
        \oc8051_xiommu1/proc_data_in [0]) ;   // aes_top.v(127)
    and (_cvpt_348, \oc8051_xiommu1/aes_top_i/n154 , \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(127)
    and (_cvpt_335, _cvpt_303, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(131)
    assign \oc8051_xiommu1/aes_top_i/aes_reg_keysel_next  = _cvpt_335 ? \oc8051_xiommu1/proc_data_in [0] : _cvpt_538;   // aes_top.v(131)
    reg2byte \oc8051_xiommu1/aes_top_i/aes_reg_opaddr_i  (.clk(clk), .rst(_cvpt_914), 
            .en(_cvpt_319), .wr(\oc8051_xiommu1/aes_top_i/n158 ), .addr(\oc8051_xiommu1/proc_addr [0]), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/aes_top_i/aes_addr_dataout }), 
            .reg_out({\oc8051_xiommu1/aes_addr }));   // aes_top.v(136)
    and (\oc8051_xiommu1/aes_top_i/n158 , _cvpt_319, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(140)
    reg2byte \oc8051_xiommu1/aes_top_i/aes_reg_oplen_i  (.clk(clk), .rst(_cvpt_914), 
            .en(_cvpt_311), .wr(\oc8051_xiommu1/aes_top_i/n159 ), .addr(\oc8051_xiommu1/proc_addr [0]), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/aes_top_i/aes_len_dataout }), 
            .reg_out({\oc8051_xiommu1/aes_len }));   // aes_top.v(150)
    and (\oc8051_xiommu1/aes_top_i/n159 , _cvpt_311, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(154)
    reg16byte \oc8051_xiommu1/aes_top_i/aes_reg_ctr_i  (.clk(clk), .rst(_cvpt_914), 
            .en(_cvpt_295), .wr(\oc8051_xiommu1/aes_top_i/n160 ), .addr({\oc8051_xiommu1/proc_addr [3:0]}), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/aes_top_i/aes_ctr_dataout }), 
            .reg_out({\oc8051_xiommu1/aes_ctr }));   // aes_top.v(167)
    and (\oc8051_xiommu1/aes_top_i/n160 , _cvpt_295, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(171)
    reg16byte \oc8051_xiommu1/aes_top_i/aes_reg_key0_i  (.clk(clk), .rst(_cvpt_914), 
            .en(_cvpt_287), .wr(\oc8051_xiommu1/aes_top_i/n161 ), .addr({\oc8051_xiommu1/proc_addr [3:0]}), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/aes_top_i/aes_key0_dataout }), 
            .reg_out({\oc8051_xiommu1/aes_key0 }));   // aes_top.v(181)
    and (\oc8051_xiommu1/aes_top_i/n161 , _cvpt_287, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(185)
    reg16byte \oc8051_xiommu1/aes_top_i/aes_reg_key1_i  (.clk(clk), .rst(_cvpt_914), 
            .en(_cvpt_279), .wr(\oc8051_xiommu1/aes_top_i/n162 ), .addr({\oc8051_xiommu1/proc_addr [3:0]}), 
            .data_in({\oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1], \oc8051_xiommu1/proc_data_in [1], 
            \oc8051_xiommu1/proc_data_in [1:0]}), .data_out({\oc8051_xiommu1/aes_top_i/aes_key1_dataout }), 
            .reg_out({\oc8051_xiommu1/aes_key1 }));   // aes_top.v(195)
    and (\oc8051_xiommu1/aes_top_i/n162 , _cvpt_279, \oc8051_xiommu1/aes_top_i/wren ) ;   // aes_top.v(199)
    and (_cvpt_336, _cvpt_530, _cvpt_402) ;   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_top_i/block_counter [4]), 
            .b(1'b1), .o(\oc8051_xiommu1/aes_top_i/n219 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n2 ));   // aes_top.v(220)
    assign \oc8051_xiommu1/aes_top_i/n178  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n165  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [15];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n179  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n166  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [14];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n180  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n167  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [13];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n181  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n168  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [12];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n182  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n169  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [11];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n183  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n170  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [10];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n184  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n171  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [9];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n185  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n172  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [8];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n186  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n173  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [7];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n187  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n174  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [6];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n188  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n175  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [5];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/n189  = _cvpt_336 ? \oc8051_xiommu1/aes_top_i/n176  : \oc8051_xiommu1/aes_top_i/operated_bytes_count [4];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [15] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n178 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [14] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n179 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [13] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n180 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [12] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n181 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [11] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n182 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [10] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n183 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [9] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n184 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [8] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n185 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [7] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n186 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [6] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n187 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [5] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n188 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [4] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n189 ;   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [3] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count [3];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [2] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count [2];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [1] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count [1];   // aes_top.v(215)
    assign \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [0] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count [0];   // aes_top.v(215)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_225/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_top_i/byte_counter [0]), 
            .b(1'b1), .o(\oc8051_xiommu1/aes_top_i/n254 ), .cout(\oc8051_xiommu1/aes_top_i/add_225/n2 ));   // aes_top.v(228)
    assign \oc8051_xiommu1/aes_top_i/n221  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n208  : \oc8051_xiommu1/aes_top_i/block_counter [15];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n222  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n209  : \oc8051_xiommu1/aes_top_i/block_counter [14];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n223  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n210  : \oc8051_xiommu1/aes_top_i/block_counter [13];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n224  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n211  : \oc8051_xiommu1/aes_top_i/block_counter [12];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n225  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n212  : \oc8051_xiommu1/aes_top_i/block_counter [11];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n226  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n213  : \oc8051_xiommu1/aes_top_i/block_counter [10];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n227  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n214  : \oc8051_xiommu1/aes_top_i/block_counter [9];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n228  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n215  : \oc8051_xiommu1/aes_top_i/block_counter [8];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n229  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n216  : \oc8051_xiommu1/aes_top_i/block_counter [7];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n230  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n217  : \oc8051_xiommu1/aes_top_i/block_counter [6];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n231  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n218  : \oc8051_xiommu1/aes_top_i/block_counter [5];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/n232  = _cvpt_364 ? \oc8051_xiommu1/aes_top_i/n219  : \oc8051_xiommu1/aes_top_i/block_counter [4];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [15] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n221 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [14] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n222 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [13] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n223 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [12] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n224 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [11] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n225 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [10] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n226 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [9] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n227 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [8] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n228 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [7] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n229 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [6] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n230 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [5] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n231 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [4] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n232 ;   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [3] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter [3];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [2] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter [2];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [1] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter [1];   // aes_top.v(221)
    assign \oc8051_xiommu1/aes_top_i/block_counter_next [0] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter [0];   // aes_top.v(221)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_240/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(231)
    assign \oc8051_xiommu1/aes_top_i/n256  = _cvpt_392 ? \oc8051_xiommu1/aes_top_i/n251  : \oc8051_xiommu1/aes_top_i/byte_counter [3];   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/n257  = _cvpt_392 ? \oc8051_xiommu1/aes_top_i/n252  : \oc8051_xiommu1/aes_top_i/byte_counter [2];   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/n258  = _cvpt_392 ? \oc8051_xiommu1/aes_top_i/n253  : \oc8051_xiommu1/aes_top_i/byte_counter [1];   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/n259  = _cvpt_392 ? \oc8051_xiommu1/aes_top_i/n254  : \oc8051_xiommu1/aes_top_i/byte_counter [0];   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/byte_counter_next [3] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n256 ;   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/byte_counter_next [2] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n257 ;   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/byte_counter_next [1] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n258 ;   // aes_top.v(229)
    assign \oc8051_xiommu1/aes_top_i/byte_counter_next [0] = _cvpt_348 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n259 ;   // aes_top.v(229)
    not (\oc8051_xiommu1/aes_top_i/n265 , \oc8051_xiommu1/aes_top_i/byte_counter [0]) ;   // aes_top.v(231)
    not (\oc8051_xiommu1/aes_top_i/n266 , \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(231)
    not (\oc8051_xiommu1/aes_top_i/n267 , \oc8051_xiommu1/aes_top_i/byte_counter [2]) ;   // aes_top.v(231)
    not (\oc8051_xiommu1/aes_top_i/n268 , \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(231)
    xor (_cvpt_3385, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [0], 
        \oc8051_xiommu1/aes_len [0]) ;   // aes_top.v(234)
    and (_cvpt_530, \oc8051_xiommu1/aes_top_i/n269 , _cvpt_392) ;   // aes_top.v(231)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_addr [0]), 
            .b(\oc8051_xiommu1/aes_top_i/block_counter [0]), .o(\oc8051_xiommu1/aes_top_i/n290 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_245/n2 ));   // aes_top.v(237)
    and (_cvpt_364, _cvpt_336, \oc8051_xiommu1/aes_top_i/n272 ) ;   // aes_top.v(234)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_top_i/n290 ), 
            .b(\oc8051_xiommu1/aes_top_i/byte_counter [0]), .o(\oc8051_xiommu1/aes_xram_addr [0]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n2 ));   // aes_top.v(237)
    or (\oc8051_xiommu1/aes_step , \oc8051_xiommu1/aes_top_i/n323 , \oc8051_xiommu1/aes_top_i/n324 ) ;   // aes_top.v(258)
    or (\oc8051_xiommu1/aes_xram_stb , _cvpt_406, _cvpt_402) ;   // aes_top.v(238)
    not (\oc8051_xiommu1/aes_top_i/aes_reg_state_next_read_data [0], _cvpt_530) ;   // aes_top.v(243)
    and (_cvpt_400, _cvpt_530, _cvpt_364) ;   // aes_top.v(247)
    assign \oc8051_xiommu1/aes_top_i/aes_reg_state_next_write_data [1] = _cvpt_400 ? 1'b0 : \oc8051_xiommu1/aes_top_i/aes_reg_state_next_read_data [0];   // aes_top.v(249)
    assign \oc8051_xiommu1/aes_top_i/aes_reg_state_next_write_data [0] = _cvpt_400 ? 1'b1 : \oc8051_xiommu1/aes_top_i/aes_reg_state_next_read_data [0];   // aes_top.v(249)
    assign \oc8051_xiommu1/aes_top_i/n315  = _cvpt_402 ? \oc8051_xiommu1/aes_top_i/aes_reg_state_next_write_data [1] : 1'b0;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/n316  = _cvpt_402 ? \oc8051_xiommu1/aes_top_i/aes_reg_state_next_write_data [0] : 1'b0;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/n317  = _cvpt_404 ? 1'b1 : \oc8051_xiommu1/aes_top_i/n315 ;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/n318  = _cvpt_404 ? 1'b1 : \oc8051_xiommu1/aes_top_i/n316 ;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/n319  = _cvpt_406 ? _cvpt_530 : \oc8051_xiommu1/aes_top_i/n317 ;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/n320  = _cvpt_406 ? \oc8051_xiommu1/aes_top_i/aes_reg_state_next_read_data [0] : \oc8051_xiommu1/aes_top_i/n318 ;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/aes_reg_state_next [1] = _cvpt_408 ? 1'b0 : \oc8051_xiommu1/aes_top_i/n319 ;   // aes_top.v(256)
    assign \oc8051_xiommu1/aes_top_i/aes_reg_state_next [0] = _cvpt_408 ? _cvpt_348 : \oc8051_xiommu1/aes_top_i/n320 ;   // aes_top.v(256)
    xor (\oc8051_xiommu1/aes_top_i/n323 , \oc8051_xiommu1/aes_state [0], 
        \oc8051_xiommu1/aes_top_i/aes_reg_state_next [0]) ;   // aes_top.v(258)
    xor (\oc8051_xiommu1/aes_top_i/n324 , \oc8051_xiommu1/aes_state [1], 
        \oc8051_xiommu1/aes_top_i/aes_reg_state_next [1]) ;   // aes_top.v(258)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_265/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(263)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_276/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(264)
    and (_cvpt_410, _cvpt_392, _cvpt_906) ;   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [7] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [7];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [6] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [6];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [5] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [5];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [4] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [4];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [3] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [3];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [2] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [2];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [1] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [1];   // aes_top.v(263)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [0] = _cvpt_410 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [0];   // aes_top.v(263)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_287/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(265)
    and (_cvpt_418, _cvpt_392, _cvpt_898) ;   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [15] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [15];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [14] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [14];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [13] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [13];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [12] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [12];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [11] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [11];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [10] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [10];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [9] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [9];   // aes_top.v(264)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [8] = _cvpt_418 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [8];   // aes_top.v(264)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_299/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(266)
    and (_cvpt_426, _cvpt_392, _cvpt_890) ;   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [23] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [23];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [22] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [22];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [21] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [21];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [20] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [20];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [19] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [19];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [18] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [18];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [17] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [17];   // aes_top.v(265)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [16] = _cvpt_426 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [16];   // aes_top.v(265)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_310/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(267)
    and (_cvpt_434, _cvpt_392, _cvpt_882) ;   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [31] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [31];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [30] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [30];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [29] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [29];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [28] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [28];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [27] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [27];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [26] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [26];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [25] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [25];   // aes_top.v(266)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [24] = _cvpt_434 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [24];   // aes_top.v(266)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_322/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(268)
    and (_cvpt_442, _cvpt_392, _cvpt_874) ;   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [39] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [39];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [38] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [38];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [37] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [37];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [36] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [36];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [35] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [35];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [34] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [34];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [33] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [33];   // aes_top.v(267)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [32] = _cvpt_442 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [32];   // aes_top.v(267)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_334/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(269)
    and (_cvpt_450, _cvpt_392, _cvpt_866) ;   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [47] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [47];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [46] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [46];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [45] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [45];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [44] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [44];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [43] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [43];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [42] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [42];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [41] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [41];   // aes_top.v(268)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [40] = _cvpt_450 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [40];   // aes_top.v(268)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_347/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(270)
    and (_cvpt_458, _cvpt_392, _cvpt_858) ;   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [55] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [55];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [54] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [54];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [53] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [53];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [52] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [52];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [51] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [51];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [50] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [50];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [49] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [49];   // aes_top.v(269)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [48] = _cvpt_458 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [48];   // aes_top.v(269)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_358/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(271)
    and (_cvpt_466, _cvpt_392, _cvpt_850) ;   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [63] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [63];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [62] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [62];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [61] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [61];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [60] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [60];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [59] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [59];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [58] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [58];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [57] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [57];   // aes_top.v(270)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [56] = _cvpt_466 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [56];   // aes_top.v(270)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_370/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(272)
    and (_cvpt_474, _cvpt_392, _cvpt_842) ;   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [71] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [71];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [70] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [70];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [69] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [69];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [68] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [68];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [67] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [67];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [66] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [66];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [65] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [65];   // aes_top.v(271)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [64] = _cvpt_474 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [64];   // aes_top.v(271)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_382/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(273)
    and (_cvpt_482, _cvpt_392, _cvpt_834) ;   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [79] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [79];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [78] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [78];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [77] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [77];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [76] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [76];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [75] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [75];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [74] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [74];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [73] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [73];   // aes_top.v(272)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [72] = _cvpt_482 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [72];   // aes_top.v(272)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_395/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(274)
    and (_cvpt_490, _cvpt_392, _cvpt_826) ;   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [87] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [87];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [86] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [86];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [85] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [85];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [84] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [84];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [83] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [83];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [82] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [82];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [81] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [81];   // aes_top.v(273)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [80] = _cvpt_490 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [80];   // aes_top.v(273)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_407/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(275)
    and (_cvpt_498, _cvpt_392, _cvpt_818) ;   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [95] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [95];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [94] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [94];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [93] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [93];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [92] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [92];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [91] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [91];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [90] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [90];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [89] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [89];   // aes_top.v(274)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [88] = _cvpt_498 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [88];   // aes_top.v(274)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_420/n1 , \oc8051_xiommu1/aes_top_i/n265 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [1]) ;   // aes_top.v(276)
    and (_cvpt_506, _cvpt_392, _cvpt_810) ;   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [103] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [103];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [102] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [102];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [101] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [101];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [100] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [100];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [99] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [99];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [98] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [98];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [97] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [97];   // aes_top.v(275)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [96] = _cvpt_506 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [96];   // aes_top.v(275)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_433/n1 , \oc8051_xiommu1/aes_top_i/byte_counter [0], 
        \oc8051_xiommu1/aes_top_i/n266 ) ;   // aes_top.v(277)
    and (_cvpt_514, _cvpt_392, _cvpt_802) ;   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [111] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [111];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [110] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [110];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [109] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [109];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [108] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [108];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [107] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [107];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [106] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [106];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [105] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [105];   // aes_top.v(276)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [104] = _cvpt_514 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [104];   // aes_top.v(276)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i1  (.cin(1'b0), .a(\oc8051_xiommu1/aes_ctr [0]), 
            .b(\oc8051_xiommu1/aes_top_i/block_counter [0]), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [0]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n2 ));   // aes_top.v(281)
    and (_cvpt_522, _cvpt_392, _cvpt_794) ;   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [119] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [119];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [118] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [118];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [117] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [117];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [116] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [116];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [115] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [115];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [114] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [114];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [113] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [113];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [112] = _cvpt_522 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [112];   // aes_top.v(277)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [127] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf [127];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [126] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf [126];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [125] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf [125];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [124] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf [124];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [123] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf [123];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [122] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf [122];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [121] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf [121];   // aes_top.v(278)
    assign \oc8051_xiommu1/aes_top_i/mem_data_buf_next [120] = _cvpt_530 ? \oc8051_xiommu1/aes_xram_data_in [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf [120];   // aes_top.v(278)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n1 , \oc8051_xiommu1/selected_port [1], 
        \oc8051_xiommu1/selected_port [2]) ;   // oc8051_memarbiter.v(126)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [0], \oc8051_xiommu1/aes_top_i/aes_out [0], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [0]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [1], \oc8051_xiommu1/aes_top_i/aes_out [1], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [1]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [2], \oc8051_xiommu1/aes_top_i/aes_out [2], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [2]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [3], \oc8051_xiommu1/aes_top_i/aes_out [3], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [3]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [4], \oc8051_xiommu1/aes_top_i/aes_out [4], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [4]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [5], \oc8051_xiommu1/aes_top_i/aes_out [5], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [5]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [6], \oc8051_xiommu1/aes_top_i/aes_out [6], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [6]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [7], \oc8051_xiommu1/aes_top_i/aes_out [7], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [7]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [8], \oc8051_xiommu1/aes_top_i/aes_out [8], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [8]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [9], \oc8051_xiommu1/aes_top_i/aes_out [9], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [9]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [10], \oc8051_xiommu1/aes_top_i/aes_out [10], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [10]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [11], \oc8051_xiommu1/aes_top_i/aes_out [11], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [11]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [12], \oc8051_xiommu1/aes_top_i/aes_out [12], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [12]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [13], \oc8051_xiommu1/aes_top_i/aes_out [13], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [13]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [14], \oc8051_xiommu1/aes_top_i/aes_out [14], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [14]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [15], \oc8051_xiommu1/aes_top_i/aes_out [15], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [15]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [16], \oc8051_xiommu1/aes_top_i/aes_out [16], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [16]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [17], \oc8051_xiommu1/aes_top_i/aes_out [17], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [17]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [18], \oc8051_xiommu1/aes_top_i/aes_out [18], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [18]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [19], \oc8051_xiommu1/aes_top_i/aes_out [19], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [19]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [20], \oc8051_xiommu1/aes_top_i/aes_out [20], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [20]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [21], \oc8051_xiommu1/aes_top_i/aes_out [21], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [21]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [22], \oc8051_xiommu1/aes_top_i/aes_out [22], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [22]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [23], \oc8051_xiommu1/aes_top_i/aes_out [23], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [23]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [24], \oc8051_xiommu1/aes_top_i/aes_out [24], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [24]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [25], \oc8051_xiommu1/aes_top_i/aes_out [25], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [25]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [26], \oc8051_xiommu1/aes_top_i/aes_out [26], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [26]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [27], \oc8051_xiommu1/aes_top_i/aes_out [27], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [27]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [28], \oc8051_xiommu1/aes_top_i/aes_out [28], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [28]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [29], \oc8051_xiommu1/aes_top_i/aes_out [29], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [29]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [30], \oc8051_xiommu1/aes_top_i/aes_out [30], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [30]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [31], \oc8051_xiommu1/aes_top_i/aes_out [31], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [31]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [32], \oc8051_xiommu1/aes_top_i/aes_out [32], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [32]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [33], \oc8051_xiommu1/aes_top_i/aes_out [33], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [33]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [34], \oc8051_xiommu1/aes_top_i/aes_out [34], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [34]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [35], \oc8051_xiommu1/aes_top_i/aes_out [35], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [35]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [36], \oc8051_xiommu1/aes_top_i/aes_out [36], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [36]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [37], \oc8051_xiommu1/aes_top_i/aes_out [37], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [37]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [38], \oc8051_xiommu1/aes_top_i/aes_out [38], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [38]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [39], \oc8051_xiommu1/aes_top_i/aes_out [39], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [39]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [40], \oc8051_xiommu1/aes_top_i/aes_out [40], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [40]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [41], \oc8051_xiommu1/aes_top_i/aes_out [41], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [41]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [42], \oc8051_xiommu1/aes_top_i/aes_out [42], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [42]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [43], \oc8051_xiommu1/aes_top_i/aes_out [43], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [43]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [44], \oc8051_xiommu1/aes_top_i/aes_out [44], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [44]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [45], \oc8051_xiommu1/aes_top_i/aes_out [45], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [45]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [46], \oc8051_xiommu1/aes_top_i/aes_out [46], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [46]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [47], \oc8051_xiommu1/aes_top_i/aes_out [47], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [47]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [48], \oc8051_xiommu1/aes_top_i/aes_out [48], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [48]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [49], \oc8051_xiommu1/aes_top_i/aes_out [49], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [49]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [50], \oc8051_xiommu1/aes_top_i/aes_out [50], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [50]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [51], \oc8051_xiommu1/aes_top_i/aes_out [51], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [51]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [52], \oc8051_xiommu1/aes_top_i/aes_out [52], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [52]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [53], \oc8051_xiommu1/aes_top_i/aes_out [53], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [53]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [54], \oc8051_xiommu1/aes_top_i/aes_out [54], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [54]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [55], \oc8051_xiommu1/aes_top_i/aes_out [55], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [55]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [56], \oc8051_xiommu1/aes_top_i/aes_out [56], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [56]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [57], \oc8051_xiommu1/aes_top_i/aes_out [57], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [57]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [58], \oc8051_xiommu1/aes_top_i/aes_out [58], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [58]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [59], \oc8051_xiommu1/aes_top_i/aes_out [59], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [59]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [60], \oc8051_xiommu1/aes_top_i/aes_out [60], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [60]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [61], \oc8051_xiommu1/aes_top_i/aes_out [61], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [61]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [62], \oc8051_xiommu1/aes_top_i/aes_out [62], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [62]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [63], \oc8051_xiommu1/aes_top_i/aes_out [63], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [63]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [64], \oc8051_xiommu1/aes_top_i/aes_out [64], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [64]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [65], \oc8051_xiommu1/aes_top_i/aes_out [65], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [65]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [66], \oc8051_xiommu1/aes_top_i/aes_out [66], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [66]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [67], \oc8051_xiommu1/aes_top_i/aes_out [67], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [67]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [68], \oc8051_xiommu1/aes_top_i/aes_out [68], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [68]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [69], \oc8051_xiommu1/aes_top_i/aes_out [69], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [69]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [70], \oc8051_xiommu1/aes_top_i/aes_out [70], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [70]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [71], \oc8051_xiommu1/aes_top_i/aes_out [71], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [71]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [72], \oc8051_xiommu1/aes_top_i/aes_out [72], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [72]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [73], \oc8051_xiommu1/aes_top_i/aes_out [73], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [73]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [74], \oc8051_xiommu1/aes_top_i/aes_out [74], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [74]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [75], \oc8051_xiommu1/aes_top_i/aes_out [75], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [75]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [76], \oc8051_xiommu1/aes_top_i/aes_out [76], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [76]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [77], \oc8051_xiommu1/aes_top_i/aes_out [77], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [77]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [78], \oc8051_xiommu1/aes_top_i/aes_out [78], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [78]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [79], \oc8051_xiommu1/aes_top_i/aes_out [79], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [79]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [80], \oc8051_xiommu1/aes_top_i/aes_out [80], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [80]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [81], \oc8051_xiommu1/aes_top_i/aes_out [81], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [81]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [82], \oc8051_xiommu1/aes_top_i/aes_out [82], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [82]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [83], \oc8051_xiommu1/aes_top_i/aes_out [83], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [83]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [84], \oc8051_xiommu1/aes_top_i/aes_out [84], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [84]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [85], \oc8051_xiommu1/aes_top_i/aes_out [85], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [85]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [86], \oc8051_xiommu1/aes_top_i/aes_out [86], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [86]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [87], \oc8051_xiommu1/aes_top_i/aes_out [87], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [87]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [88], \oc8051_xiommu1/aes_top_i/aes_out [88], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [88]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [89], \oc8051_xiommu1/aes_top_i/aes_out [89], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [89]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [90], \oc8051_xiommu1/aes_top_i/aes_out [90], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [90]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [91], \oc8051_xiommu1/aes_top_i/aes_out [91], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [91]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [92], \oc8051_xiommu1/aes_top_i/aes_out [92], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [92]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [93], \oc8051_xiommu1/aes_top_i/aes_out [93], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [93]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [94], \oc8051_xiommu1/aes_top_i/aes_out [94], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [94]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [95], \oc8051_xiommu1/aes_top_i/aes_out [95], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [95]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [96], \oc8051_xiommu1/aes_top_i/aes_out [96], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [96]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [97], \oc8051_xiommu1/aes_top_i/aes_out [97], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [97]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [98], \oc8051_xiommu1/aes_top_i/aes_out [98], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [98]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [99], \oc8051_xiommu1/aes_top_i/aes_out [99], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [99]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [100], \oc8051_xiommu1/aes_top_i/aes_out [100], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [100]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [101], \oc8051_xiommu1/aes_top_i/aes_out [101], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [101]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [102], \oc8051_xiommu1/aes_top_i/aes_out [102], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [102]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [103], \oc8051_xiommu1/aes_top_i/aes_out [103], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [103]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [104], \oc8051_xiommu1/aes_top_i/aes_out [104], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [104]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [105], \oc8051_xiommu1/aes_top_i/aes_out [105], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [105]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [106], \oc8051_xiommu1/aes_top_i/aes_out [106], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [106]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [107], \oc8051_xiommu1/aes_top_i/aes_out [107], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [107]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [108], \oc8051_xiommu1/aes_top_i/aes_out [108], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [108]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [109], \oc8051_xiommu1/aes_top_i/aes_out [109], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [109]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [110], \oc8051_xiommu1/aes_top_i/aes_out [110], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [110]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [111], \oc8051_xiommu1/aes_top_i/aes_out [111], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [111]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [112], \oc8051_xiommu1/aes_top_i/aes_out [112], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [112]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [113], \oc8051_xiommu1/aes_top_i/aes_out [113], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [113]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [114], \oc8051_xiommu1/aes_top_i/aes_out [114], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [114]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [115], \oc8051_xiommu1/aes_top_i/aes_out [115], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [115]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [116], \oc8051_xiommu1/aes_top_i/aes_out [116], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [116]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [117], \oc8051_xiommu1/aes_top_i/aes_out [117], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [117]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [118], \oc8051_xiommu1/aes_top_i/aes_out [118], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [118]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [119], \oc8051_xiommu1/aes_top_i/aes_out [119], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [119]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [120], \oc8051_xiommu1/aes_top_i/aes_out [120], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [120]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [121], \oc8051_xiommu1/aes_top_i/aes_out [121], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [121]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [122], \oc8051_xiommu1/aes_top_i/aes_out [122], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [122]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [123], \oc8051_xiommu1/aes_top_i/aes_out [123], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [123]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [124], \oc8051_xiommu1/aes_top_i/aes_out [124], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [124]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [125], \oc8051_xiommu1/aes_top_i/aes_out [125], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [125]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [126], \oc8051_xiommu1/aes_top_i/aes_out [126], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [126]) ;   // aes_top.v(283)
    xor (\oc8051_xiommu1/aes_top_i/encrypted_data [127], \oc8051_xiommu1/aes_top_i/aes_out [127], 
        \oc8051_xiommu1/aes_top_i/mem_data_buf [127]) ;   // aes_top.v(283)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [127] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [127] : \oc8051_xiommu1/aes_key0 [127];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [126] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [126] : \oc8051_xiommu1/aes_key0 [126];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [125] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [125] : \oc8051_xiommu1/aes_key0 [125];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [124] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [124] : \oc8051_xiommu1/aes_key0 [124];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [123] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [123] : \oc8051_xiommu1/aes_key0 [123];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [122] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [122] : \oc8051_xiommu1/aes_key0 [122];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [121] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [121] : \oc8051_xiommu1/aes_key0 [121];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [120] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [120] : \oc8051_xiommu1/aes_key0 [120];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [119] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [119] : \oc8051_xiommu1/aes_key0 [119];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [118] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [118] : \oc8051_xiommu1/aes_key0 [118];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [117] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [117] : \oc8051_xiommu1/aes_key0 [117];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [116] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [116] : \oc8051_xiommu1/aes_key0 [116];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [115] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [115] : \oc8051_xiommu1/aes_key0 [115];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [114] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [114] : \oc8051_xiommu1/aes_key0 [114];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [113] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [113] : \oc8051_xiommu1/aes_key0 [113];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [112] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [112] : \oc8051_xiommu1/aes_key0 [112];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [111] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [111] : \oc8051_xiommu1/aes_key0 [111];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [110] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [110] : \oc8051_xiommu1/aes_key0 [110];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [109] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [109] : \oc8051_xiommu1/aes_key0 [109];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [108] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [108] : \oc8051_xiommu1/aes_key0 [108];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [107] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [107] : \oc8051_xiommu1/aes_key0 [107];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [106] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [106] : \oc8051_xiommu1/aes_key0 [106];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [105] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [105] : \oc8051_xiommu1/aes_key0 [105];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [104] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [104] : \oc8051_xiommu1/aes_key0 [104];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [103] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [103] : \oc8051_xiommu1/aes_key0 [103];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [102] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [102] : \oc8051_xiommu1/aes_key0 [102];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [101] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [101] : \oc8051_xiommu1/aes_key0 [101];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [100] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [100] : \oc8051_xiommu1/aes_key0 [100];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [99] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [99] : \oc8051_xiommu1/aes_key0 [99];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [98] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [98] : \oc8051_xiommu1/aes_key0 [98];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [97] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [97] : \oc8051_xiommu1/aes_key0 [97];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [96] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [96] : \oc8051_xiommu1/aes_key0 [96];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [95] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [95] : \oc8051_xiommu1/aes_key0 [95];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [94] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [94] : \oc8051_xiommu1/aes_key0 [94];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [93] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [93] : \oc8051_xiommu1/aes_key0 [93];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [92] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [92] : \oc8051_xiommu1/aes_key0 [92];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [91] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [91] : \oc8051_xiommu1/aes_key0 [91];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [90] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [90] : \oc8051_xiommu1/aes_key0 [90];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [89] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [89] : \oc8051_xiommu1/aes_key0 [89];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [88] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [88] : \oc8051_xiommu1/aes_key0 [88];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [87] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [87] : \oc8051_xiommu1/aes_key0 [87];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [86] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [86] : \oc8051_xiommu1/aes_key0 [86];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [85] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [85] : \oc8051_xiommu1/aes_key0 [85];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [84] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [84] : \oc8051_xiommu1/aes_key0 [84];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [83] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [83] : \oc8051_xiommu1/aes_key0 [83];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [82] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [82] : \oc8051_xiommu1/aes_key0 [82];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [81] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [81] : \oc8051_xiommu1/aes_key0 [81];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [80] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [80] : \oc8051_xiommu1/aes_key0 [80];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [79] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [79] : \oc8051_xiommu1/aes_key0 [79];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [78] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [78] : \oc8051_xiommu1/aes_key0 [78];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [77] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [77] : \oc8051_xiommu1/aes_key0 [77];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [76] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [76] : \oc8051_xiommu1/aes_key0 [76];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [75] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [75] : \oc8051_xiommu1/aes_key0 [75];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [74] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [74] : \oc8051_xiommu1/aes_key0 [74];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [73] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [73] : \oc8051_xiommu1/aes_key0 [73];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [72] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [72] : \oc8051_xiommu1/aes_key0 [72];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [71] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [71] : \oc8051_xiommu1/aes_key0 [71];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [70] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [70] : \oc8051_xiommu1/aes_key0 [70];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [69] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [69] : \oc8051_xiommu1/aes_key0 [69];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [68] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [68] : \oc8051_xiommu1/aes_key0 [68];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [67] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [67] : \oc8051_xiommu1/aes_key0 [67];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [66] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [66] : \oc8051_xiommu1/aes_key0 [66];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [65] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [65] : \oc8051_xiommu1/aes_key0 [65];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [64] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [64] : \oc8051_xiommu1/aes_key0 [64];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [63] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [63] : \oc8051_xiommu1/aes_key0 [63];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [62] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [62] : \oc8051_xiommu1/aes_key0 [62];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [61] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [61] : \oc8051_xiommu1/aes_key0 [61];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [60] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [60] : \oc8051_xiommu1/aes_key0 [60];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [59] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [59] : \oc8051_xiommu1/aes_key0 [59];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [58] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [58] : \oc8051_xiommu1/aes_key0 [58];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [57] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [57] : \oc8051_xiommu1/aes_key0 [57];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [56] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [56] : \oc8051_xiommu1/aes_key0 [56];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [55] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [55] : \oc8051_xiommu1/aes_key0 [55];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [54] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [54] : \oc8051_xiommu1/aes_key0 [54];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [53] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [53] : \oc8051_xiommu1/aes_key0 [53];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [52] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [52] : \oc8051_xiommu1/aes_key0 [52];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [51] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [51] : \oc8051_xiommu1/aes_key0 [51];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [50] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [50] : \oc8051_xiommu1/aes_key0 [50];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [49] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [49] : \oc8051_xiommu1/aes_key0 [49];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [48] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [48] : \oc8051_xiommu1/aes_key0 [48];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [47] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [47] : \oc8051_xiommu1/aes_key0 [47];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [46] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [46] : \oc8051_xiommu1/aes_key0 [46];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [45] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [45] : \oc8051_xiommu1/aes_key0 [45];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [44] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [44] : \oc8051_xiommu1/aes_key0 [44];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [43] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [43] : \oc8051_xiommu1/aes_key0 [43];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [42] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [42] : \oc8051_xiommu1/aes_key0 [42];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [41] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [41] : \oc8051_xiommu1/aes_key0 [41];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [40] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [40] : \oc8051_xiommu1/aes_key0 [40];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [39] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [39] : \oc8051_xiommu1/aes_key0 [39];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [38] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [38] : \oc8051_xiommu1/aes_key0 [38];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [37] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [37] : \oc8051_xiommu1/aes_key0 [37];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [36] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [36] : \oc8051_xiommu1/aes_key0 [36];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [35] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [35] : \oc8051_xiommu1/aes_key0 [35];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [34] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [34] : \oc8051_xiommu1/aes_key0 [34];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [33] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [33] : \oc8051_xiommu1/aes_key0 [33];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [32] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [32] : \oc8051_xiommu1/aes_key0 [32];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [31] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [31] : \oc8051_xiommu1/aes_key0 [31];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [30] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [30] : \oc8051_xiommu1/aes_key0 [30];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [29] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [29] : \oc8051_xiommu1/aes_key0 [29];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [28] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [28] : \oc8051_xiommu1/aes_key0 [28];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [27] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [27] : \oc8051_xiommu1/aes_key0 [27];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [26] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [26] : \oc8051_xiommu1/aes_key0 [26];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [25] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [25] : \oc8051_xiommu1/aes_key0 [25];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [24] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [24] : \oc8051_xiommu1/aes_key0 [24];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [23] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [23] : \oc8051_xiommu1/aes_key0 [23];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [22] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [22] : \oc8051_xiommu1/aes_key0 [22];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [21] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [21] : \oc8051_xiommu1/aes_key0 [21];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [20] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [20] : \oc8051_xiommu1/aes_key0 [20];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [19] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [19] : \oc8051_xiommu1/aes_key0 [19];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [18] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [18] : \oc8051_xiommu1/aes_key0 [18];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [17] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [17] : \oc8051_xiommu1/aes_key0 [17];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [16] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [16] : \oc8051_xiommu1/aes_key0 [16];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [15] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [15] : \oc8051_xiommu1/aes_key0 [15];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [14] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [14] : \oc8051_xiommu1/aes_key0 [14];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [13] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [13] : \oc8051_xiommu1/aes_key0 [13];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [12] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [12] : \oc8051_xiommu1/aes_key0 [12];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [11] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [11] : \oc8051_xiommu1/aes_key0 [11];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [10] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [10] : \oc8051_xiommu1/aes_key0 [10];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [9] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [9] : \oc8051_xiommu1/aes_key0 [9];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [8] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [8] : \oc8051_xiommu1/aes_key0 [8];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [7] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [7] : \oc8051_xiommu1/aes_key0 [7];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [6] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [6] : \oc8051_xiommu1/aes_key0 [6];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [5] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [5] : \oc8051_xiommu1/aes_key0 [5];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [4] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [4] : \oc8051_xiommu1/aes_key0 [4];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [3] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [3] : \oc8051_xiommu1/aes_key0 [3];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [2] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [2] : \oc8051_xiommu1/aes_key0 [2];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [1] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [1] : \oc8051_xiommu1/aes_key0 [1];   // aes_top.v(284)
    assign \oc8051_xiommu1/aes_top_i/aes_curr_key [0] = _cvpt_538 ? \oc8051_xiommu1/aes_key1 [0] : \oc8051_xiommu1/aes_key0 [0];   // aes_top.v(284)
    aes_128 \oc8051_xiommu1/aes_top_i/aes_128_i  (.clk(clk), .state({\oc8051_xiommu1/aes_top_i/aes_ctr_v }), 
            .key({\oc8051_xiommu1/aes_top_i/aes_curr_key }), .out({\oc8051_xiommu1/aes_top_i/aes_out }));   // aes_top.v(285)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [127] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [127] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [127];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [126] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [126] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [126];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [125] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [125] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [125];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [124] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [124] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [124];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [123] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [123] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [123];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [122] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [122] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [122];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [121] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [121] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [121];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [120] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [120] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [120];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [119] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [119] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [119];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [118] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [118] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [118];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [117] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [117] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [117];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [116] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [116] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [116];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [115] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [115] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [115];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [114] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [114] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [114];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [113] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [113] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [113];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [112] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [112] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [112];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [111] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [111] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [111];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [110] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [110] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [110];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [109] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [109] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [109];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [108] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [108] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [108];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [107] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [107] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [107];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [106] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [106] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [106];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [105] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [105] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [105];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [104] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [104] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [104];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [103] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [103] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [103];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [102] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [102] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [102];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [101] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [101] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [101];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [100] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [100] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [100];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [99] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [99] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [99];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [98] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [98] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [98];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [97] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [97] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [97];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [96] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [96] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [96];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [95] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [95] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [95];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [94] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [94] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [94];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [93] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [93] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [93];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [92] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [92] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [92];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [91] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [91] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [91];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [90] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [90] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [90];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [89] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [89] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [89];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [88] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [88] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [88];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [87] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [87] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [87];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [86] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [86] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [86];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [85] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [85] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [85];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [84] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [84] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [84];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [83] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [83] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [83];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [82] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [82] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [82];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [81] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [81] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [81];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [80] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [80] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [80];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [79] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [79] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [79];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [78] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [78] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [78];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [77] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [77] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [77];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [76] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [76] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [76];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [75] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [75] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [75];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [74] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [74] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [74];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [73] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [73] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [73];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [72] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [72] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [72];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [71] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [71] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [71];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [70] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [70] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [70];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [69] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [69] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [69];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [68] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [68] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [68];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [67] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [67] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [67];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [66] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [66] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [66];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [65] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [65] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [65];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [64] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [64] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [64];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [63] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [63] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [63];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [62] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [62] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [62];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [61] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [61] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [61];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [60] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [60] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [60];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [59] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [59] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [59];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [58] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [58] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [58];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [57] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [57] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [57];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [56] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [56] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [56];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [55] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [55] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [55];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [54] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [54] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [54];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [53] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [53] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [53];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [52] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [52] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [52];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [51] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [51] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [51];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [50] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [50] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [50];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [49] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [49] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [49];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [48] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [48] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [48];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [47] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [47] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [47];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [46] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [46] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [46];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [45] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [45] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [45];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [44] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [44] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [44];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [43] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [43] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [43];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [42] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [42] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [42];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [41] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [41] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [41];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [40] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [40] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [40];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [39] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [39] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [39];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [38] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [38] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [38];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [37] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [37] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [37];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [36] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [36] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [36];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [35] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [35] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [35];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [34] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [34] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [34];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [33] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [33] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [33];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [32] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [32] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [32];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [31] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [31] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [31];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [30] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [30] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [30];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [29] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [29] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [29];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [28] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [28] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [28];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [27] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [27] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [27];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [26] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [26] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [26];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [25] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [25] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [25];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [24] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [24] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [24];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [23] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [23] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [23];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [22] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [22] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [22];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [21] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [21] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [21];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [20] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [20] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [20];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [19] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [19] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [19];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [18] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [18] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [18];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [17] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [17] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [17];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [16] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [16] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [16];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [15] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [15] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [15];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [14] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [14] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [14];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [13] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [13] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [13];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [12] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [12] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [12];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [11] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [11] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [11];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [10] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [10] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [10];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [9] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [9] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [9];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [8] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [8] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [8];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [7] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [7] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [7];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [6] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [6] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [6];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [5] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [5] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [5];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [4] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [4] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [4];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [3] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [3] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [3];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [2] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [2] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [2];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [1] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [1] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [1];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [0] = _cvpt_404 ? \oc8051_xiommu1/aes_top_i/encrypted_data [0] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [0];   // aes_top.v(296)
    assign \oc8051_xiommu1/aes_top_i/n1074  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [119] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [127];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1075  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [118] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [126];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1076  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [117] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [125];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1077  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [116] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [124];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1078  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [115] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [123];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1079  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [114] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [122];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1080  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [113] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [121];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1081  = _cvpt_794 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [112] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf [120];   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1082  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [111] : \oc8051_xiommu1/aes_top_i/n1074 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1083  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [110] : \oc8051_xiommu1/aes_top_i/n1075 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1084  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [109] : \oc8051_xiommu1/aes_top_i/n1076 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1085  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [108] : \oc8051_xiommu1/aes_top_i/n1077 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1086  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [107] : \oc8051_xiommu1/aes_top_i/n1078 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1087  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [106] : \oc8051_xiommu1/aes_top_i/n1079 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1088  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [105] : \oc8051_xiommu1/aes_top_i/n1080 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1089  = _cvpt_802 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [104] : \oc8051_xiommu1/aes_top_i/n1081 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1090  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [103] : \oc8051_xiommu1/aes_top_i/n1082 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1091  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [102] : \oc8051_xiommu1/aes_top_i/n1083 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1092  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [101] : \oc8051_xiommu1/aes_top_i/n1084 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1093  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [100] : \oc8051_xiommu1/aes_top_i/n1085 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1094  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [99] : \oc8051_xiommu1/aes_top_i/n1086 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1095  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [98] : \oc8051_xiommu1/aes_top_i/n1087 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1096  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [97] : \oc8051_xiommu1/aes_top_i/n1088 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1097  = _cvpt_810 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [96] : \oc8051_xiommu1/aes_top_i/n1089 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1098  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [95] : \oc8051_xiommu1/aes_top_i/n1090 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1099  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [94] : \oc8051_xiommu1/aes_top_i/n1091 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1100  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [93] : \oc8051_xiommu1/aes_top_i/n1092 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1101  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [92] : \oc8051_xiommu1/aes_top_i/n1093 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1102  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [91] : \oc8051_xiommu1/aes_top_i/n1094 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1103  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [90] : \oc8051_xiommu1/aes_top_i/n1095 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1104  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [89] : \oc8051_xiommu1/aes_top_i/n1096 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1105  = _cvpt_818 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [88] : \oc8051_xiommu1/aes_top_i/n1097 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1106  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [87] : \oc8051_xiommu1/aes_top_i/n1098 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1107  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [86] : \oc8051_xiommu1/aes_top_i/n1099 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1108  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [85] : \oc8051_xiommu1/aes_top_i/n1100 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1109  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [84] : \oc8051_xiommu1/aes_top_i/n1101 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1110  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [83] : \oc8051_xiommu1/aes_top_i/n1102 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1111  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [82] : \oc8051_xiommu1/aes_top_i/n1103 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1112  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [81] : \oc8051_xiommu1/aes_top_i/n1104 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1113  = _cvpt_826 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [80] : \oc8051_xiommu1/aes_top_i/n1105 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1114  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [79] : \oc8051_xiommu1/aes_top_i/n1106 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1115  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [78] : \oc8051_xiommu1/aes_top_i/n1107 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1116  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [77] : \oc8051_xiommu1/aes_top_i/n1108 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1117  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [76] : \oc8051_xiommu1/aes_top_i/n1109 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1118  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [75] : \oc8051_xiommu1/aes_top_i/n1110 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1119  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [74] : \oc8051_xiommu1/aes_top_i/n1111 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1120  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [73] : \oc8051_xiommu1/aes_top_i/n1112 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1121  = _cvpt_834 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [72] : \oc8051_xiommu1/aes_top_i/n1113 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1122  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [71] : \oc8051_xiommu1/aes_top_i/n1114 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1123  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [70] : \oc8051_xiommu1/aes_top_i/n1115 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1124  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [69] : \oc8051_xiommu1/aes_top_i/n1116 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1125  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [68] : \oc8051_xiommu1/aes_top_i/n1117 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1126  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [67] : \oc8051_xiommu1/aes_top_i/n1118 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1127  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [66] : \oc8051_xiommu1/aes_top_i/n1119 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1128  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [65] : \oc8051_xiommu1/aes_top_i/n1120 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1129  = _cvpt_842 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [64] : \oc8051_xiommu1/aes_top_i/n1121 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1130  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [63] : \oc8051_xiommu1/aes_top_i/n1122 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1131  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [62] : \oc8051_xiommu1/aes_top_i/n1123 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1132  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [61] : \oc8051_xiommu1/aes_top_i/n1124 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1133  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [60] : \oc8051_xiommu1/aes_top_i/n1125 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1134  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [59] : \oc8051_xiommu1/aes_top_i/n1126 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1135  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [58] : \oc8051_xiommu1/aes_top_i/n1127 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1136  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [57] : \oc8051_xiommu1/aes_top_i/n1128 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1137  = _cvpt_850 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [56] : \oc8051_xiommu1/aes_top_i/n1129 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1138  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [55] : \oc8051_xiommu1/aes_top_i/n1130 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1139  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [54] : \oc8051_xiommu1/aes_top_i/n1131 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1140  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [53] : \oc8051_xiommu1/aes_top_i/n1132 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1141  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [52] : \oc8051_xiommu1/aes_top_i/n1133 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1142  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [51] : \oc8051_xiommu1/aes_top_i/n1134 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1143  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [50] : \oc8051_xiommu1/aes_top_i/n1135 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1144  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [49] : \oc8051_xiommu1/aes_top_i/n1136 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1145  = _cvpt_858 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [48] : \oc8051_xiommu1/aes_top_i/n1137 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1146  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [47] : \oc8051_xiommu1/aes_top_i/n1138 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1147  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [46] : \oc8051_xiommu1/aes_top_i/n1139 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1148  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [45] : \oc8051_xiommu1/aes_top_i/n1140 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1149  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [44] : \oc8051_xiommu1/aes_top_i/n1141 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1150  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [43] : \oc8051_xiommu1/aes_top_i/n1142 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1151  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [42] : \oc8051_xiommu1/aes_top_i/n1143 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1152  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [41] : \oc8051_xiommu1/aes_top_i/n1144 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1153  = _cvpt_866 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [40] : \oc8051_xiommu1/aes_top_i/n1145 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1154  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [39] : \oc8051_xiommu1/aes_top_i/n1146 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1155  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [38] : \oc8051_xiommu1/aes_top_i/n1147 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1156  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [37] : \oc8051_xiommu1/aes_top_i/n1148 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1157  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [36] : \oc8051_xiommu1/aes_top_i/n1149 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1158  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [35] : \oc8051_xiommu1/aes_top_i/n1150 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1159  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [34] : \oc8051_xiommu1/aes_top_i/n1151 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1160  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [33] : \oc8051_xiommu1/aes_top_i/n1152 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1161  = _cvpt_874 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [32] : \oc8051_xiommu1/aes_top_i/n1153 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1162  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [31] : \oc8051_xiommu1/aes_top_i/n1154 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1163  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [30] : \oc8051_xiommu1/aes_top_i/n1155 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1164  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [29] : \oc8051_xiommu1/aes_top_i/n1156 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1165  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [28] : \oc8051_xiommu1/aes_top_i/n1157 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1166  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [27] : \oc8051_xiommu1/aes_top_i/n1158 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1167  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [26] : \oc8051_xiommu1/aes_top_i/n1159 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1168  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [25] : \oc8051_xiommu1/aes_top_i/n1160 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1169  = _cvpt_882 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [24] : \oc8051_xiommu1/aes_top_i/n1161 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1170  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [23] : \oc8051_xiommu1/aes_top_i/n1162 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1171  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [22] : \oc8051_xiommu1/aes_top_i/n1163 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1172  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [21] : \oc8051_xiommu1/aes_top_i/n1164 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1173  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [20] : \oc8051_xiommu1/aes_top_i/n1165 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1174  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [19] : \oc8051_xiommu1/aes_top_i/n1166 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1175  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [18] : \oc8051_xiommu1/aes_top_i/n1167 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1176  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [17] : \oc8051_xiommu1/aes_top_i/n1168 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1177  = _cvpt_890 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [16] : \oc8051_xiommu1/aes_top_i/n1169 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1178  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [15] : \oc8051_xiommu1/aes_top_i/n1170 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1179  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [14] : \oc8051_xiommu1/aes_top_i/n1171 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1180  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [13] : \oc8051_xiommu1/aes_top_i/n1172 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1181  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [12] : \oc8051_xiommu1/aes_top_i/n1173 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1182  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [11] : \oc8051_xiommu1/aes_top_i/n1174 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1183  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [10] : \oc8051_xiommu1/aes_top_i/n1175 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1184  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [9] : \oc8051_xiommu1/aes_top_i/n1176 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1185  = _cvpt_898 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [8] : \oc8051_xiommu1/aes_top_i/n1177 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [7] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [7] : \oc8051_xiommu1/aes_top_i/n1178 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [6] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [6] : \oc8051_xiommu1/aes_top_i/n1179 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [5] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [5] : \oc8051_xiommu1/aes_top_i/n1180 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [4] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [4] : \oc8051_xiommu1/aes_top_i/n1181 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [3] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [3] : \oc8051_xiommu1/aes_top_i/n1182 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [2] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [2] : \oc8051_xiommu1/aes_top_i/n1183 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [1] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [1] : \oc8051_xiommu1/aes_top_i/n1184 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_xram_data_out [0] = _cvpt_906 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [0] : \oc8051_xiommu1/aes_top_i/n1185 ;   // aes_top.v(314)
    assign \oc8051_xiommu1/aes_top_i/n1195  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/aes_reg_state_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1196  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/aes_reg_state_next [0];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1197  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [15];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1198  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [14];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1199  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [13];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1200  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [12];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1201  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [11];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1202  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [10];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1203  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [9];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1204  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [8];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1205  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [7];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1206  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [6];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1207  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [5];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1208  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [4];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1209  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [3];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1210  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [2];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1211  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1212  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/block_counter_next [0];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1213  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/byte_counter_next [3];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1214  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/byte_counter_next [2];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1215  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/byte_counter_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1216  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/byte_counter_next [0];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1217  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [15];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1218  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [14];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1219  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [13];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1220  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [12];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1221  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [11];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1222  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [10];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1223  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [9];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1224  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [8];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1225  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [7];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1226  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [6];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1227  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [5];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1228  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [4];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1229  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [3];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1230  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [2];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1231  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1232  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [0];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1233  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/aes_top_i/aes_reg_keysel_next ;   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1234  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [127] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [127];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1235  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [126] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [126];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1236  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [125] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [125];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1237  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [124] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [124];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1238  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [123] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [123];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1239  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [122] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [122];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1240  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [121] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [121];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1241  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [120] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [120];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1242  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [119] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [119];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1243  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [118] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [118];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1244  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [117] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [117];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1245  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [116] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [116];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1246  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [115] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [115];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1247  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [114] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [114];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1248  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [113] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [113];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1249  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [112] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [112];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1250  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [111] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [111];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1251  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [110] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [110];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1252  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [109] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [109];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1253  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [108] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [108];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1254  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [107] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [107];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1255  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [106] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [106];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1256  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [105] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [105];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1257  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [104] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [104];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1258  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [103] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [103];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1259  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [102] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [102];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1260  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [101] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [101];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1261  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [100] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [100];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1262  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [99] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [99];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1263  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [98] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [98];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1264  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [97] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [97];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1265  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [96] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [96];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1266  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [95] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [95];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1267  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [94] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [94];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1268  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [93] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [93];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1269  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [92] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [92];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1270  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [91] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [91];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1271  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [90] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [90];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1272  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [89] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [89];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1273  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [88] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [88];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1274  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [87] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [87];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1275  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [86] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [86];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1276  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [85] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [85];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1277  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [84] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [84];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1278  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [83] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [83];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1279  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [82] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [82];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1280  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [81] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [81];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1281  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [80] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [80];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1282  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [79] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [79];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1283  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [78] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [78];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1284  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [77] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [77];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1285  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [76] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [76];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1286  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [75] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [75];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1287  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [74] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [74];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1288  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [73] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [73];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1289  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [72] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [72];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1290  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [71] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [71];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1291  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [70] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [70];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1292  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [69] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [69];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1293  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [68] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [68];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1294  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [67] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [67];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1295  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [66] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [66];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1296  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [65] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [65];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1297  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [64] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [64];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1298  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [63] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [63];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1299  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [62] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [62];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1300  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [61] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [61];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1301  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [60] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [60];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1302  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [59] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [59];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1303  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [58] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [58];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1304  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [57] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [57];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1305  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [56] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [56];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1306  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [55] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [55];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1307  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [54] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [54];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1308  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [53] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [53];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1309  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [52] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [52];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1310  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [51] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [51];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1311  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [50] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [50];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1312  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [49] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [49];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1313  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [48] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [48];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1314  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [47] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [47];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1315  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [46] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [46];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1316  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [45] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [45];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1317  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [44] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [44];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1318  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [43] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [43];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1319  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [42] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [42];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1320  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [41] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [41];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1321  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [40] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [40];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1322  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [39] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [39];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1323  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [38] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [38];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1324  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [37] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [37];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1325  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [36] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [36];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1326  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [35] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [35];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1327  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [34] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [34];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1328  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [33] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [33];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1329  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [32] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [32];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1330  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [31] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [31];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1331  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [30] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [30];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1332  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [29] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [29];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1333  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [28] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [28];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1334  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [27] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [27];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1335  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [26] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [26];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1336  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [25] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [25];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1337  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [24] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [24];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1338  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [23] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [23];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1339  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [22] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [22];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1340  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [21] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [21];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1341  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [20] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [20];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1342  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [19] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [19];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1343  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [18] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [18];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1344  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [17] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [17];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1345  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [16] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [16];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1346  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [15] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [15];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1347  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [14] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [14];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1348  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [13] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [13];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1349  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [12] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [12];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1350  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [11] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [11];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1351  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [10] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [10];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1352  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [9] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [9];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1353  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [8] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [8];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1354  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [7] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [7];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1355  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [6] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [6];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1356  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [5] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [5];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1357  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [4] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [4];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1358  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [3] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [3];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1359  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [2] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [2];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1360  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [1] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1361  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/mem_data_buf [0] : \oc8051_xiommu1/aes_top_i/mem_data_buf_next [0];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1362  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [127] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [127];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1363  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [126] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [126];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1364  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [125] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [125];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1365  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [124] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [124];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1366  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [123] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [123];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1367  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [122] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [122];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1368  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [121] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [121];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1369  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [120] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [120];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1370  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [119] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [119];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1371  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [118] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [118];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1372  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [117] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [117];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1373  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [116] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [116];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1374  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [115] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [115];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1375  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [114] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [114];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1376  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [113] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [113];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1377  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [112] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [112];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1378  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [111] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [111];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1379  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [110] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [110];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1380  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [109] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [109];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1381  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [108] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [108];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1382  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [107] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [107];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1383  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [106] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [106];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1384  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [105] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [105];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1385  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [104] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [104];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1386  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [103] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [103];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1387  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [102] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [102];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1388  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [101] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [101];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1389  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [100] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [100];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1390  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [99] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [99];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1391  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [98] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [98];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1392  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [97] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [97];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1393  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [96] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [96];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1394  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [95] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [95];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1395  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [94] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [94];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1396  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [93] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [93];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1397  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [92] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [92];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1398  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [91] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [91];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1399  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [90] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [90];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1400  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [89] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [89];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1401  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [88] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [88];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1402  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [87] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [87];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1403  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [86] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [86];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1404  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [85] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [85];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1405  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [84] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [84];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1406  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [83] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [83];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1407  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [82] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [82];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1408  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [81] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [81];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1409  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [80] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [80];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1410  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [79] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [79];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1411  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [78] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [78];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1412  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [77] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [77];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1413  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [76] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [76];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1414  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [75] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [75];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1415  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [74] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [74];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1416  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [73] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [73];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1417  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [72] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [72];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1418  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [71] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [71];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1419  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [70] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [70];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1420  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [69] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [69];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1421  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [68] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [68];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1422  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [67] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [67];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1423  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [66] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [66];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1424  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [65] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [65];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1425  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [64] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [64];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1426  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [63] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [63];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1427  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [62] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [62];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1428  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [61] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [61];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1429  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [60] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [60];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1430  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [59] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [59];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1431  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [58] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [58];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1432  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [57] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [57];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1433  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [56] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [56];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1434  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [55] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [55];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1435  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [54] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [54];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1436  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [53] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [53];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1437  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [52] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [52];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1438  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [51] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [51];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1439  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [50] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [50];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1440  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [49] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [49];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1441  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [48] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [48];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1442  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [47] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [47];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1443  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [46] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [46];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1444  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [45] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [45];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1445  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [44] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [44];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1446  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [43] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [43];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1447  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [42] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [42];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1448  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [41] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [41];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1449  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [40] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [40];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1450  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [39] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [39];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1451  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [38] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [38];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1452  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [37] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [37];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1453  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [36] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [36];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1454  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [35] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [35];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1455  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [34] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [34];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1456  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [33] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [33];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1457  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [32] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [32];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1458  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [31] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [31];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1459  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [30] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [30];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1460  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [29] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [29];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1461  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [28] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [28];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1462  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [27] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [27];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1463  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [26] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [26];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1464  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [25] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [25];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1465  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [24] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [24];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1466  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [23] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [23];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1467  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [22] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [22];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1468  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [21] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [21];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1469  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [20] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [20];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1470  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [19] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [19];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1471  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [18] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [18];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1472  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [17] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [17];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1473  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [16] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [16];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1474  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [15] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [15];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1475  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [14] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [14];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1476  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [13] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [13];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1477  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [12] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [12];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1478  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [11] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [11];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1479  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [10] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [10];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1480  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [9] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [9];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1481  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [8] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [8];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1482  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [7] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [7];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1483  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [6] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [6];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1484  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [5] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [5];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1485  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [4] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [4];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1486  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [3] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [3];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1487  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [2] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [2];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1488  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [1] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [1];   // aes_top.v(335)
    assign \oc8051_xiommu1/aes_top_i/n1489  = _cvpt_914 ? \oc8051_xiommu1/aes_top_i/encrypted_data_buf [0] : \oc8051_xiommu1/aes_top_i/encrypted_data_buf_next [0];   // aes_top.v(335)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1303  (.d(\oc8051_xiommu1/aes_top_i/n1196 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_state [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1304  (.d(\oc8051_xiommu1/aes_top_i/n1197 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [15]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1305  (.d(\oc8051_xiommu1/aes_top_i/n1198 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [14]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1306  (.d(\oc8051_xiommu1/aes_top_i/n1199 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [13]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1307  (.d(\oc8051_xiommu1/aes_top_i/n1200 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [12]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1308  (.d(\oc8051_xiommu1/aes_top_i/n1201 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [11]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1309  (.d(\oc8051_xiommu1/aes_top_i/n1202 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [10]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1310  (.d(\oc8051_xiommu1/aes_top_i/n1203 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [9]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1311  (.d(\oc8051_xiommu1/aes_top_i/n1204 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [8]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1312  (.d(\oc8051_xiommu1/aes_top_i/n1205 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [7]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1313  (.d(\oc8051_xiommu1/aes_top_i/n1206 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [6]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1314  (.d(\oc8051_xiommu1/aes_top_i/n1207 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [5]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1315  (.d(\oc8051_xiommu1/aes_top_i/n1208 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [4]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1316  (.d(\oc8051_xiommu1/aes_top_i/n1209 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [3]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1317  (.d(\oc8051_xiommu1/aes_top_i/n1210 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [2]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1318  (.d(\oc8051_xiommu1/aes_top_i/n1211 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [1]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1319  (.d(\oc8051_xiommu1/aes_top_i/n1212 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/block_counter [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1320  (.d(\oc8051_xiommu1/aes_top_i/n1213 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/byte_counter [3]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1321  (.d(\oc8051_xiommu1/aes_top_i/n1214 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/byte_counter [2]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1322  (.d(\oc8051_xiommu1/aes_top_i/n1215 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/byte_counter [1]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1323  (.d(\oc8051_xiommu1/aes_top_i/n1216 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/byte_counter [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1324  (.d(\oc8051_xiommu1/aes_top_i/n1217 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [15]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1325  (.d(\oc8051_xiommu1/aes_top_i/n1218 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [14]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1326  (.d(\oc8051_xiommu1/aes_top_i/n1219 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [13]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1327  (.d(\oc8051_xiommu1/aes_top_i/n1220 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [12]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1328  (.d(\oc8051_xiommu1/aes_top_i/n1221 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [11]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1329  (.d(\oc8051_xiommu1/aes_top_i/n1222 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [10]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1330  (.d(\oc8051_xiommu1/aes_top_i/n1223 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [9]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1331  (.d(\oc8051_xiommu1/aes_top_i/n1224 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [8]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1332  (.d(\oc8051_xiommu1/aes_top_i/n1225 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [7]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1333  (.d(\oc8051_xiommu1/aes_top_i/n1226 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [6]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1334  (.d(\oc8051_xiommu1/aes_top_i/n1227 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [5]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1335  (.d(\oc8051_xiommu1/aes_top_i/n1228 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [4]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1336  (.d(\oc8051_xiommu1/aes_top_i/n1229 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [3]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1337  (.d(\oc8051_xiommu1/aes_top_i/n1230 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [2]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1338  (.d(\oc8051_xiommu1/aes_top_i/n1231 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [1]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1339  (.d(\oc8051_xiommu1/aes_top_i/n1232 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/operated_bytes_count [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1340  (.d(\oc8051_xiommu1/aes_top_i/n1233 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(_cvpt_538));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1341  (.d(\oc8051_xiommu1/aes_top_i/n1234 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [127]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1342  (.d(\oc8051_xiommu1/aes_top_i/n1235 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [126]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1343  (.d(\oc8051_xiommu1/aes_top_i/n1236 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [125]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1344  (.d(\oc8051_xiommu1/aes_top_i/n1237 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [124]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1345  (.d(\oc8051_xiommu1/aes_top_i/n1238 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [123]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1346  (.d(\oc8051_xiommu1/aes_top_i/n1239 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [122]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1347  (.d(\oc8051_xiommu1/aes_top_i/n1240 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [121]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1348  (.d(\oc8051_xiommu1/aes_top_i/n1241 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [120]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1349  (.d(\oc8051_xiommu1/aes_top_i/n1242 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [119]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1350  (.d(\oc8051_xiommu1/aes_top_i/n1243 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [118]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1351  (.d(\oc8051_xiommu1/aes_top_i/n1244 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [117]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1352  (.d(\oc8051_xiommu1/aes_top_i/n1245 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [116]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1353  (.d(\oc8051_xiommu1/aes_top_i/n1246 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [115]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1354  (.d(\oc8051_xiommu1/aes_top_i/n1247 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [114]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1355  (.d(\oc8051_xiommu1/aes_top_i/n1248 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [113]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1356  (.d(\oc8051_xiommu1/aes_top_i/n1249 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [112]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1357  (.d(\oc8051_xiommu1/aes_top_i/n1250 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [111]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1358  (.d(\oc8051_xiommu1/aes_top_i/n1251 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [110]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1359  (.d(\oc8051_xiommu1/aes_top_i/n1252 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [109]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1360  (.d(\oc8051_xiommu1/aes_top_i/n1253 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [108]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1361  (.d(\oc8051_xiommu1/aes_top_i/n1254 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [107]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1362  (.d(\oc8051_xiommu1/aes_top_i/n1255 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [106]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1363  (.d(\oc8051_xiommu1/aes_top_i/n1256 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [105]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1364  (.d(\oc8051_xiommu1/aes_top_i/n1257 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [104]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1365  (.d(\oc8051_xiommu1/aes_top_i/n1258 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [103]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1366  (.d(\oc8051_xiommu1/aes_top_i/n1259 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [102]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1367  (.d(\oc8051_xiommu1/aes_top_i/n1260 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [101]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1368  (.d(\oc8051_xiommu1/aes_top_i/n1261 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [100]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1369  (.d(\oc8051_xiommu1/aes_top_i/n1262 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [99]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1370  (.d(\oc8051_xiommu1/aes_top_i/n1263 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [98]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1371  (.d(\oc8051_xiommu1/aes_top_i/n1264 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [97]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1372  (.d(\oc8051_xiommu1/aes_top_i/n1265 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [96]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1373  (.d(\oc8051_xiommu1/aes_top_i/n1266 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [95]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1374  (.d(\oc8051_xiommu1/aes_top_i/n1267 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [94]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1375  (.d(\oc8051_xiommu1/aes_top_i/n1268 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [93]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1376  (.d(\oc8051_xiommu1/aes_top_i/n1269 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [92]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1377  (.d(\oc8051_xiommu1/aes_top_i/n1270 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [91]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1378  (.d(\oc8051_xiommu1/aes_top_i/n1271 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [90]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1379  (.d(\oc8051_xiommu1/aes_top_i/n1272 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [89]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1380  (.d(\oc8051_xiommu1/aes_top_i/n1273 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [88]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1381  (.d(\oc8051_xiommu1/aes_top_i/n1274 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [87]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1382  (.d(\oc8051_xiommu1/aes_top_i/n1275 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [86]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1383  (.d(\oc8051_xiommu1/aes_top_i/n1276 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [85]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1384  (.d(\oc8051_xiommu1/aes_top_i/n1277 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [84]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1385  (.d(\oc8051_xiommu1/aes_top_i/n1278 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [83]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1386  (.d(\oc8051_xiommu1/aes_top_i/n1279 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [82]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1387  (.d(\oc8051_xiommu1/aes_top_i/n1280 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [81]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1388  (.d(\oc8051_xiommu1/aes_top_i/n1281 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [80]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1389  (.d(\oc8051_xiommu1/aes_top_i/n1282 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [79]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1390  (.d(\oc8051_xiommu1/aes_top_i/n1283 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [78]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1391  (.d(\oc8051_xiommu1/aes_top_i/n1284 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [77]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1392  (.d(\oc8051_xiommu1/aes_top_i/n1285 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [76]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1393  (.d(\oc8051_xiommu1/aes_top_i/n1286 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [75]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1394  (.d(\oc8051_xiommu1/aes_top_i/n1287 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [74]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1395  (.d(\oc8051_xiommu1/aes_top_i/n1288 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [73]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1396  (.d(\oc8051_xiommu1/aes_top_i/n1289 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [72]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1397  (.d(\oc8051_xiommu1/aes_top_i/n1290 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [71]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1398  (.d(\oc8051_xiommu1/aes_top_i/n1291 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [70]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1399  (.d(\oc8051_xiommu1/aes_top_i/n1292 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [69]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1400  (.d(\oc8051_xiommu1/aes_top_i/n1293 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [68]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1401  (.d(\oc8051_xiommu1/aes_top_i/n1294 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [67]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1402  (.d(\oc8051_xiommu1/aes_top_i/n1295 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [66]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1403  (.d(\oc8051_xiommu1/aes_top_i/n1296 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [65]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1404  (.d(\oc8051_xiommu1/aes_top_i/n1297 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [64]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1405  (.d(\oc8051_xiommu1/aes_top_i/n1298 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [63]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1406  (.d(\oc8051_xiommu1/aes_top_i/n1299 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [62]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1407  (.d(\oc8051_xiommu1/aes_top_i/n1300 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [61]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1408  (.d(\oc8051_xiommu1/aes_top_i/n1301 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [60]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1409  (.d(\oc8051_xiommu1/aes_top_i/n1302 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [59]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1410  (.d(\oc8051_xiommu1/aes_top_i/n1303 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [58]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1411  (.d(\oc8051_xiommu1/aes_top_i/n1304 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [57]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1412  (.d(\oc8051_xiommu1/aes_top_i/n1305 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [56]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1413  (.d(\oc8051_xiommu1/aes_top_i/n1306 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [55]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1414  (.d(\oc8051_xiommu1/aes_top_i/n1307 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [54]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1415  (.d(\oc8051_xiommu1/aes_top_i/n1308 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [53]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1416  (.d(\oc8051_xiommu1/aes_top_i/n1309 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [52]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1417  (.d(\oc8051_xiommu1/aes_top_i/n1310 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [51]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1418  (.d(\oc8051_xiommu1/aes_top_i/n1311 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [50]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1419  (.d(\oc8051_xiommu1/aes_top_i/n1312 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [49]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1420  (.d(\oc8051_xiommu1/aes_top_i/n1313 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [48]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1421  (.d(\oc8051_xiommu1/aes_top_i/n1314 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [47]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1422  (.d(\oc8051_xiommu1/aes_top_i/n1315 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [46]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1423  (.d(\oc8051_xiommu1/aes_top_i/n1316 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [45]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1424  (.d(\oc8051_xiommu1/aes_top_i/n1317 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [44]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1425  (.d(\oc8051_xiommu1/aes_top_i/n1318 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [43]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1426  (.d(\oc8051_xiommu1/aes_top_i/n1319 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [42]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1427  (.d(\oc8051_xiommu1/aes_top_i/n1320 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [41]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1428  (.d(\oc8051_xiommu1/aes_top_i/n1321 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [40]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1429  (.d(\oc8051_xiommu1/aes_top_i/n1322 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [39]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1430  (.d(\oc8051_xiommu1/aes_top_i/n1323 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [38]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1431  (.d(\oc8051_xiommu1/aes_top_i/n1324 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [37]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1432  (.d(\oc8051_xiommu1/aes_top_i/n1325 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [36]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1433  (.d(\oc8051_xiommu1/aes_top_i/n1326 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [35]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1434  (.d(\oc8051_xiommu1/aes_top_i/n1327 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [34]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1435  (.d(\oc8051_xiommu1/aes_top_i/n1328 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [33]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1436  (.d(\oc8051_xiommu1/aes_top_i/n1329 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [32]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1437  (.d(\oc8051_xiommu1/aes_top_i/n1330 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [31]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1438  (.d(\oc8051_xiommu1/aes_top_i/n1331 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [30]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1439  (.d(\oc8051_xiommu1/aes_top_i/n1332 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [29]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1440  (.d(\oc8051_xiommu1/aes_top_i/n1333 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [28]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1441  (.d(\oc8051_xiommu1/aes_top_i/n1334 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [27]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1442  (.d(\oc8051_xiommu1/aes_top_i/n1335 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [26]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1443  (.d(\oc8051_xiommu1/aes_top_i/n1336 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [25]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1444  (.d(\oc8051_xiommu1/aes_top_i/n1337 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [24]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1445  (.d(\oc8051_xiommu1/aes_top_i/n1338 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [23]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1446  (.d(\oc8051_xiommu1/aes_top_i/n1339 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [22]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1447  (.d(\oc8051_xiommu1/aes_top_i/n1340 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [21]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1448  (.d(\oc8051_xiommu1/aes_top_i/n1341 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [20]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1449  (.d(\oc8051_xiommu1/aes_top_i/n1342 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [19]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1450  (.d(\oc8051_xiommu1/aes_top_i/n1343 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [18]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1451  (.d(\oc8051_xiommu1/aes_top_i/n1344 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [17]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1452  (.d(\oc8051_xiommu1/aes_top_i/n1345 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [16]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1453  (.d(\oc8051_xiommu1/aes_top_i/n1346 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [15]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1454  (.d(\oc8051_xiommu1/aes_top_i/n1347 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [14]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1455  (.d(\oc8051_xiommu1/aes_top_i/n1348 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [13]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1456  (.d(\oc8051_xiommu1/aes_top_i/n1349 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [12]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1457  (.d(\oc8051_xiommu1/aes_top_i/n1350 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [11]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1458  (.d(\oc8051_xiommu1/aes_top_i/n1351 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [10]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1459  (.d(\oc8051_xiommu1/aes_top_i/n1352 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [9]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1460  (.d(\oc8051_xiommu1/aes_top_i/n1353 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [8]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1461  (.d(\oc8051_xiommu1/aes_top_i/n1354 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [7]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1462  (.d(\oc8051_xiommu1/aes_top_i/n1355 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [6]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1463  (.d(\oc8051_xiommu1/aes_top_i/n1356 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [5]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1464  (.d(\oc8051_xiommu1/aes_top_i/n1357 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [4]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1465  (.d(\oc8051_xiommu1/aes_top_i/n1358 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [3]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1466  (.d(\oc8051_xiommu1/aes_top_i/n1359 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [2]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1467  (.d(\oc8051_xiommu1/aes_top_i/n1360 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [1]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1468  (.d(\oc8051_xiommu1/aes_top_i/n1361 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/mem_data_buf [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1469  (.d(\oc8051_xiommu1/aes_top_i/n1362 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [127]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1470  (.d(\oc8051_xiommu1/aes_top_i/n1363 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [126]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1471  (.d(\oc8051_xiommu1/aes_top_i/n1364 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [125]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1472  (.d(\oc8051_xiommu1/aes_top_i/n1365 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [124]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1473  (.d(\oc8051_xiommu1/aes_top_i/n1366 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [123]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1474  (.d(\oc8051_xiommu1/aes_top_i/n1367 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [122]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1475  (.d(\oc8051_xiommu1/aes_top_i/n1368 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [121]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1476  (.d(\oc8051_xiommu1/aes_top_i/n1369 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [120]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1477  (.d(\oc8051_xiommu1/aes_top_i/n1370 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [119]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1478  (.d(\oc8051_xiommu1/aes_top_i/n1371 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [118]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1479  (.d(\oc8051_xiommu1/aes_top_i/n1372 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [117]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1480  (.d(\oc8051_xiommu1/aes_top_i/n1373 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [116]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1481  (.d(\oc8051_xiommu1/aes_top_i/n1374 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [115]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1482  (.d(\oc8051_xiommu1/aes_top_i/n1375 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [114]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1483  (.d(\oc8051_xiommu1/aes_top_i/n1376 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [113]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1484  (.d(\oc8051_xiommu1/aes_top_i/n1377 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [112]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1485  (.d(\oc8051_xiommu1/aes_top_i/n1378 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [111]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1486  (.d(\oc8051_xiommu1/aes_top_i/n1379 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [110]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1487  (.d(\oc8051_xiommu1/aes_top_i/n1380 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [109]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1488  (.d(\oc8051_xiommu1/aes_top_i/n1381 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [108]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1489  (.d(\oc8051_xiommu1/aes_top_i/n1382 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [107]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1490  (.d(\oc8051_xiommu1/aes_top_i/n1383 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [106]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1491  (.d(\oc8051_xiommu1/aes_top_i/n1384 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [105]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1492  (.d(\oc8051_xiommu1/aes_top_i/n1385 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [104]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1493  (.d(\oc8051_xiommu1/aes_top_i/n1386 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [103]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1494  (.d(\oc8051_xiommu1/aes_top_i/n1387 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [102]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1495  (.d(\oc8051_xiommu1/aes_top_i/n1388 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [101]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1496  (.d(\oc8051_xiommu1/aes_top_i/n1389 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [100]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1497  (.d(\oc8051_xiommu1/aes_top_i/n1390 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [99]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1498  (.d(\oc8051_xiommu1/aes_top_i/n1391 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [98]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1499  (.d(\oc8051_xiommu1/aes_top_i/n1392 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [97]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1500  (.d(\oc8051_xiommu1/aes_top_i/n1393 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [96]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1501  (.d(\oc8051_xiommu1/aes_top_i/n1394 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [95]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1502  (.d(\oc8051_xiommu1/aes_top_i/n1395 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [94]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1503  (.d(\oc8051_xiommu1/aes_top_i/n1396 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [93]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1504  (.d(\oc8051_xiommu1/aes_top_i/n1397 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [92]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1505  (.d(\oc8051_xiommu1/aes_top_i/n1398 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [91]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1506  (.d(\oc8051_xiommu1/aes_top_i/n1399 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [90]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1507  (.d(\oc8051_xiommu1/aes_top_i/n1400 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [89]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1508  (.d(\oc8051_xiommu1/aes_top_i/n1401 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [88]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1509  (.d(\oc8051_xiommu1/aes_top_i/n1402 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [87]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1510  (.d(\oc8051_xiommu1/aes_top_i/n1403 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [86]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1511  (.d(\oc8051_xiommu1/aes_top_i/n1404 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [85]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1512  (.d(\oc8051_xiommu1/aes_top_i/n1405 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [84]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1513  (.d(\oc8051_xiommu1/aes_top_i/n1406 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [83]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1514  (.d(\oc8051_xiommu1/aes_top_i/n1407 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [82]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1515  (.d(\oc8051_xiommu1/aes_top_i/n1408 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [81]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1516  (.d(\oc8051_xiommu1/aes_top_i/n1409 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [80]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1517  (.d(\oc8051_xiommu1/aes_top_i/n1410 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [79]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1518  (.d(\oc8051_xiommu1/aes_top_i/n1411 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [78]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1519  (.d(\oc8051_xiommu1/aes_top_i/n1412 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [77]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1520  (.d(\oc8051_xiommu1/aes_top_i/n1413 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [76]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1521  (.d(\oc8051_xiommu1/aes_top_i/n1414 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [75]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1522  (.d(\oc8051_xiommu1/aes_top_i/n1415 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [74]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1523  (.d(\oc8051_xiommu1/aes_top_i/n1416 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [73]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1524  (.d(\oc8051_xiommu1/aes_top_i/n1417 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [72]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1525  (.d(\oc8051_xiommu1/aes_top_i/n1418 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [71]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1526  (.d(\oc8051_xiommu1/aes_top_i/n1419 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [70]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1527  (.d(\oc8051_xiommu1/aes_top_i/n1420 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [69]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1528  (.d(\oc8051_xiommu1/aes_top_i/n1421 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [68]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1529  (.d(\oc8051_xiommu1/aes_top_i/n1422 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [67]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1530  (.d(\oc8051_xiommu1/aes_top_i/n1423 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [66]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1531  (.d(\oc8051_xiommu1/aes_top_i/n1424 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [65]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1532  (.d(\oc8051_xiommu1/aes_top_i/n1425 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [64]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1533  (.d(\oc8051_xiommu1/aes_top_i/n1426 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [63]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1534  (.d(\oc8051_xiommu1/aes_top_i/n1427 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [62]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1535  (.d(\oc8051_xiommu1/aes_top_i/n1428 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [61]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1536  (.d(\oc8051_xiommu1/aes_top_i/n1429 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [60]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1537  (.d(\oc8051_xiommu1/aes_top_i/n1430 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [59]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1538  (.d(\oc8051_xiommu1/aes_top_i/n1431 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [58]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1539  (.d(\oc8051_xiommu1/aes_top_i/n1432 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [57]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1540  (.d(\oc8051_xiommu1/aes_top_i/n1433 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [56]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1541  (.d(\oc8051_xiommu1/aes_top_i/n1434 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [55]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1542  (.d(\oc8051_xiommu1/aes_top_i/n1435 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [54]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1543  (.d(\oc8051_xiommu1/aes_top_i/n1436 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [53]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1544  (.d(\oc8051_xiommu1/aes_top_i/n1437 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [52]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1545  (.d(\oc8051_xiommu1/aes_top_i/n1438 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [51]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1546  (.d(\oc8051_xiommu1/aes_top_i/n1439 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [50]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1547  (.d(\oc8051_xiommu1/aes_top_i/n1440 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [49]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1548  (.d(\oc8051_xiommu1/aes_top_i/n1441 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [48]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1549  (.d(\oc8051_xiommu1/aes_top_i/n1442 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [47]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1550  (.d(\oc8051_xiommu1/aes_top_i/n1443 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [46]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1551  (.d(\oc8051_xiommu1/aes_top_i/n1444 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [45]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1552  (.d(\oc8051_xiommu1/aes_top_i/n1445 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [44]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1553  (.d(\oc8051_xiommu1/aes_top_i/n1446 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [43]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1554  (.d(\oc8051_xiommu1/aes_top_i/n1447 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [42]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1555  (.d(\oc8051_xiommu1/aes_top_i/n1448 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [41]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1556  (.d(\oc8051_xiommu1/aes_top_i/n1449 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [40]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1557  (.d(\oc8051_xiommu1/aes_top_i/n1450 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [39]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1558  (.d(\oc8051_xiommu1/aes_top_i/n1451 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [38]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1559  (.d(\oc8051_xiommu1/aes_top_i/n1452 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [37]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1560  (.d(\oc8051_xiommu1/aes_top_i/n1453 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [36]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1561  (.d(\oc8051_xiommu1/aes_top_i/n1454 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [35]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1562  (.d(\oc8051_xiommu1/aes_top_i/n1455 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [34]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1563  (.d(\oc8051_xiommu1/aes_top_i/n1456 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [33]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1564  (.d(\oc8051_xiommu1/aes_top_i/n1457 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [32]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1565  (.d(\oc8051_xiommu1/aes_top_i/n1458 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [31]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1566  (.d(\oc8051_xiommu1/aes_top_i/n1459 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [30]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1567  (.d(\oc8051_xiommu1/aes_top_i/n1460 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [29]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1568  (.d(\oc8051_xiommu1/aes_top_i/n1461 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [28]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1569  (.d(\oc8051_xiommu1/aes_top_i/n1462 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [27]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1570  (.d(\oc8051_xiommu1/aes_top_i/n1463 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [26]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1571  (.d(\oc8051_xiommu1/aes_top_i/n1464 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [25]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1572  (.d(\oc8051_xiommu1/aes_top_i/n1465 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [24]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1573  (.d(\oc8051_xiommu1/aes_top_i/n1466 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [23]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1574  (.d(\oc8051_xiommu1/aes_top_i/n1467 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [22]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1575  (.d(\oc8051_xiommu1/aes_top_i/n1468 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [21]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1576  (.d(\oc8051_xiommu1/aes_top_i/n1469 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [20]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1577  (.d(\oc8051_xiommu1/aes_top_i/n1470 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [19]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1578  (.d(\oc8051_xiommu1/aes_top_i/n1471 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [18]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1579  (.d(\oc8051_xiommu1/aes_top_i/n1472 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [17]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1580  (.d(\oc8051_xiommu1/aes_top_i/n1473 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [16]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1581  (.d(\oc8051_xiommu1/aes_top_i/n1474 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [15]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1582  (.d(\oc8051_xiommu1/aes_top_i/n1475 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [14]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1583  (.d(\oc8051_xiommu1/aes_top_i/n1476 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [13]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1584  (.d(\oc8051_xiommu1/aes_top_i/n1477 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [12]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1585  (.d(\oc8051_xiommu1/aes_top_i/n1478 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [11]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1586  (.d(\oc8051_xiommu1/aes_top_i/n1479 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [10]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1587  (.d(\oc8051_xiommu1/aes_top_i/n1480 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [9]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1588  (.d(\oc8051_xiommu1/aes_top_i/n1481 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [8]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1589  (.d(\oc8051_xiommu1/aes_top_i/n1482 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [7]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1590  (.d(\oc8051_xiommu1/aes_top_i/n1483 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [6]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1591  (.d(\oc8051_xiommu1/aes_top_i/n1484 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [5]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1592  (.d(\oc8051_xiommu1/aes_top_i/n1485 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [4]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1593  (.d(\oc8051_xiommu1/aes_top_i/n1486 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [3]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1594  (.d(\oc8051_xiommu1/aes_top_i/n1487 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [2]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1595  (.d(\oc8051_xiommu1/aes_top_i/n1488 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [1]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1596  (.d(\oc8051_xiommu1/aes_top_i/n1489 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_top_i/encrypted_data_buf [0]));   // aes_top.v(336)
    VERIFIC_DFFRS \oc8051_xiommu1/aes_top_i/i1302  (.d(\oc8051_xiommu1/aes_top_i/n1195 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/aes_state [1]));   // aes_top.v(336)
    assign \oc8051_xiommu1/proc_stb  = _cvpt_1209 ? \oc8051_xiommu1/proc1_stb_xram  : \oc8051_xiommu1/proc0_stb_xram ;   // oc8051_procarbiter.v(89)
    assign \oc8051_xiommu1/proc_wr  = _cvpt_1209 ? \oc8051_xiommu1/write1_xram  : \oc8051_xiommu1/write0_xram ;   // oc8051_procarbiter.v(91)
    assign \oc8051_xiommu1/proc_addr [15] = _cvpt_1209 ? ext_addr[15] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [14] = _cvpt_1209 ? ext_addr[14] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [13] = _cvpt_1209 ? ext_addr[13] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [12] = _cvpt_1209 ? ext_addr[12] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [11] = _cvpt_1209 ? ext_addr[11] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [10] = _cvpt_1209 ? ext_addr[10] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [9] = _cvpt_1209 ? ext_addr[9] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [8] = _cvpt_1209 ? ext_addr[8] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [7] = _cvpt_1209 ? ext_addr[7] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [6] = _cvpt_1209 ? ext_addr[6] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [5] = _cvpt_1209 ? ext_addr[5] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [4] = _cvpt_1209 ? ext_addr[4] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [3] = _cvpt_1209 ? ext_addr[3] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [2] = _cvpt_1209 ? ext_addr[2] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [1] = _cvpt_1209 ? ext_addr[1] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_addr [0] = _cvpt_1209 ? ext_addr[0] : p3_in[2];   // oc8051_procarbiter.v(93)
    assign \oc8051_xiommu1/proc_data_in [0] = _cvpt_1209 ? data_out[0] : p3_in[2];   // oc8051_procarbiter.v(95)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/ack_A  = _cvpt_1209 ? \oc8051_xiommu1/proc_ack  : 1'b0;   // oc8051_procarbiter.v(97)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/ack_B  = _cvpt_1209 ? 1'b0 : \oc8051_xiommu1/proc_ack ;   // oc8051_procarbiter.v(98)
    assign \oc8051_xiommu1/priv_lvl  = _cvpt_1209 ? p3_in[2] : priv_lvl;   // oc8051_procarbiter.v(103)
    assign \oc8051_xiommu1/dpc_ot [15] = _cvpt_1209 ? p3_in[2] : dpc_ot[15];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [14] = _cvpt_1209 ? p3_in[2] : dpc_ot[14];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [13] = _cvpt_1209 ? p3_in[2] : dpc_ot[13];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [12] = _cvpt_1209 ? p3_in[2] : dpc_ot[12];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [11] = _cvpt_1209 ? p3_in[2] : dpc_ot[11];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [10] = _cvpt_1209 ? p3_in[2] : dpc_ot[10];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [9] = _cvpt_1209 ? p3_in[2] : dpc_ot[9];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [8] = _cvpt_1209 ? p3_in[2] : dpc_ot[8];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [7] = _cvpt_1209 ? p3_in[2] : dpc_ot[7];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [6] = _cvpt_1209 ? p3_in[2] : dpc_ot[6];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [5] = _cvpt_1209 ? p3_in[2] : dpc_ot[5];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [4] = _cvpt_1209 ? p3_in[2] : dpc_ot[4];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [3] = _cvpt_1209 ? p3_in[2] : dpc_ot[3];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [2] = _cvpt_1209 ? p3_in[2] : dpc_ot[2];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [1] = _cvpt_1209 ? p3_in[2] : dpc_ot[1];   // oc8051_procarbiter.v(105)
    assign \oc8051_xiommu1/dpc_ot [0] = _cvpt_1209 ? p3_in[2] : dpc_ot[0];   // oc8051_procarbiter.v(105)
    not (\oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_inuse_next , \oc8051_xiommu1/proc_ack ) ;   // oc8051_procarbiter.v(111)
    or (\oc8051_xiommu1/oc8051_procarbiter_i/n58 , \oc8051_xiommu1/proc1_stb_xram , 
        \oc8051_xiommu1/proc0_stb_xram ) ;   // oc8051_procarbiter.v(115)
    and (\oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_idle_next , \oc8051_xiommu1/oc8051_procarbiter_i/n58 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_inuse_next ) ;   // oc8051_procarbiter.v(115)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_next  = _cvpt_1247 ? \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_inuse_next  : \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_idle_next ;   // oc8051_procarbiter.v(120)
    not (\oc8051_xiommu1/oc8051_procarbiter_i/n64 , _cvpt_1247) ;   // oc8051_procarbiter.v(123)
    and (_cvpt_1248, \oc8051_xiommu1/oc8051_procarbiter_i/n64 , \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_next ) ;   // oc8051_procarbiter.v(123)
    and (\oc8051_xiommu1/oc8051_procarbiter_i/n67 , \oc8051_xiommu1/proc1_stb_xram , 
        \oc8051_xiommu1/proc0_stb_xram ) ;   // oc8051_procarbiter.v(128)
    and (\oc8051_xiommu1/oc8051_procarbiter_i/n69 , \oc8051_xiommu1/oc8051_procarbiter_i/n67 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder ) ;   // oc8051_procarbiter.v(128)
    not (\oc8051_xiommu1/oc8051_procarbiter_i/n70 , \oc8051_xiommu1/proc1_stb_xram ) ;   // oc8051_procarbiter.v(128)
    and (\oc8051_xiommu1/oc8051_procarbiter_i/n71 , \oc8051_xiommu1/oc8051_procarbiter_i/n70 , 
        \oc8051_xiommu1/proc0_stb_xram ) ;   // oc8051_procarbiter.v(128)
    or (\oc8051_xiommu1/oc8051_procarbiter_i/n72 , \oc8051_xiommu1/oc8051_procarbiter_i/n69 , 
        \oc8051_xiommu1/oc8051_procarbiter_i/n71 ) ;   // oc8051_procarbiter.v(128)
    not (\oc8051_xiommu1/oc8051_procarbiter_i/arbit_winner , \oc8051_xiommu1/oc8051_procarbiter_i/n72 ) ;   // oc8051_procarbiter.v(128)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder_next  = _cvpt_1248 ? \oc8051_xiommu1/oc8051_procarbiter_i/arbit_winner  : \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder ;   // oc8051_procarbiter.v(138)
    assign _cvpt_1209 = _cvpt_1247 ? \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder  : \oc8051_xiommu1/oc8051_procarbiter_i/arbit_winner ;   // oc8051_procarbiter.v(142)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/n78  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_procarbiter_i/arbiter_state_next ;   // oc8051_procarbiter.v(154)
    assign \oc8051_xiommu1/oc8051_procarbiter_i/n79  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder_next ;   // oc8051_procarbiter.v(154)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_procarbiter_i/i81  (.d(\oc8051_xiommu1/oc8051_procarbiter_i/n79 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_procarbiter_i/arbit_holder ));   // oc8051_procarbiter.v(155)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_procarbiter_i/i80  (.d(\oc8051_xiommu1/oc8051_procarbiter_i/n78 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(_cvpt_1247));   // oc8051_procarbiter.v(155)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n1 , \oc8051_xiommu1/selected_port [1], 
        \oc8051_xiommu1/selected_port [2]) ;   // oc8051_memarbiter.v(127)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n5 , \oc8051_xiommu1/selected_port [0]) ;   // oc8051_memarbiter.v(127)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/n7 , 
        \oc8051_xiommu1/selected_port [2]) ;   // oc8051_memarbiter.v(128)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n7 , \oc8051_xiommu1/selected_port [1]) ;   // oc8051_memarbiter.v(128)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n1 , \oc8051_xiommu1/oc8051_memarbiter_i/n7 , 
        \oc8051_xiommu1/selected_port [2]) ;   // oc8051_memarbiter.v(129)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n1 , \oc8051_xiommu1/selected_port [1], 
        \oc8051_xiommu1/oc8051_memarbiter_i/n152 ) ;   // oc8051_memarbiter.v(150)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n12  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_stb  : \oc8051_xiommu1/memwr_xram_stb ;   // oc8051_memarbiter.v(129)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n13  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_stb  : \oc8051_xiommu1/oc8051_memarbiter_i/n12 ;   // oc8051_memarbiter.v(129)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n14  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_stb  : \oc8051_xiommu1/oc8051_memarbiter_i/n13 ;   // oc8051_memarbiter.v(129)
    assign \oc8051_xiommu1/stb_out  = _cvpt_1255 ? \oc8051_xiommu1/proc_stb  : \oc8051_xiommu1/oc8051_memarbiter_i/n14 ;   // oc8051_memarbiter.v(129)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n24  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_wr  : \oc8051_xiommu1/memwr_xram_wr ;   // oc8051_memarbiter.v(134)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n25  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_wr  : \oc8051_xiommu1/oc8051_memarbiter_i/n24 ;   // oc8051_memarbiter.v(134)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n26  = _cvpt_1254 ? _cvpt_402 : \oc8051_xiommu1/oc8051_memarbiter_i/n25 ;   // oc8051_memarbiter.v(134)
    assign \oc8051_xiommu1/wr_out  = _cvpt_1255 ? \oc8051_xiommu1/proc_wr  : \oc8051_xiommu1/oc8051_memarbiter_i/n26 ;   // oc8051_memarbiter.v(134)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n36  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [15] : \oc8051_xiommu1/memwr_xram_addr [15];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n37  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [14] : \oc8051_xiommu1/memwr_xram_addr [14];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n38  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [13] : \oc8051_xiommu1/memwr_xram_addr [13];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n39  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [12] : \oc8051_xiommu1/memwr_xram_addr [12];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n40  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [11] : \oc8051_xiommu1/memwr_xram_addr [11];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n41  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [10] : \oc8051_xiommu1/memwr_xram_addr [10];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n42  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [9] : \oc8051_xiommu1/memwr_xram_addr [9];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n43  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [8] : \oc8051_xiommu1/memwr_xram_addr [8];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n44  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [7] : \oc8051_xiommu1/memwr_xram_addr [7];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n45  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [6] : \oc8051_xiommu1/memwr_xram_addr [6];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n46  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [5] : \oc8051_xiommu1/memwr_xram_addr [5];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n47  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [4] : \oc8051_xiommu1/memwr_xram_addr [4];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n48  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [3] : \oc8051_xiommu1/memwr_xram_addr [3];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n49  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [2] : \oc8051_xiommu1/memwr_xram_addr [2];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n50  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [1] : \oc8051_xiommu1/memwr_xram_addr [1];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n51  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_addr [0] : \oc8051_xiommu1/memwr_xram_addr [0];   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n52  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [15] : \oc8051_xiommu1/oc8051_memarbiter_i/n36 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n53  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [14] : \oc8051_xiommu1/oc8051_memarbiter_i/n37 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n54  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [13] : \oc8051_xiommu1/oc8051_memarbiter_i/n38 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n55  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [12] : \oc8051_xiommu1/oc8051_memarbiter_i/n39 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n56  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [11] : \oc8051_xiommu1/oc8051_memarbiter_i/n40 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n57  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [10] : \oc8051_xiommu1/oc8051_memarbiter_i/n41 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n58  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [9] : \oc8051_xiommu1/oc8051_memarbiter_i/n42 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n59  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [8] : \oc8051_xiommu1/oc8051_memarbiter_i/n43 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n60  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [7] : \oc8051_xiommu1/oc8051_memarbiter_i/n44 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n61  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [6] : \oc8051_xiommu1/oc8051_memarbiter_i/n45 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n62  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [5] : \oc8051_xiommu1/oc8051_memarbiter_i/n46 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n63  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [4] : \oc8051_xiommu1/oc8051_memarbiter_i/n47 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n64  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [3] : \oc8051_xiommu1/oc8051_memarbiter_i/n48 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n65  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [2] : \oc8051_xiommu1/oc8051_memarbiter_i/n49 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n66  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n50 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n67  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_addr [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n51 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n68  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [15] : \oc8051_xiommu1/oc8051_memarbiter_i/n52 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n69  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [14] : \oc8051_xiommu1/oc8051_memarbiter_i/n53 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n70  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [13] : \oc8051_xiommu1/oc8051_memarbiter_i/n54 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n71  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [12] : \oc8051_xiommu1/oc8051_memarbiter_i/n55 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n72  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [11] : \oc8051_xiommu1/oc8051_memarbiter_i/n56 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n73  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [10] : \oc8051_xiommu1/oc8051_memarbiter_i/n57 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n74  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [9] : \oc8051_xiommu1/oc8051_memarbiter_i/n58 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n75  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [8] : \oc8051_xiommu1/oc8051_memarbiter_i/n59 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n76  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [7] : \oc8051_xiommu1/oc8051_memarbiter_i/n60 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n77  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [6] : \oc8051_xiommu1/oc8051_memarbiter_i/n61 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n78  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [5] : \oc8051_xiommu1/oc8051_memarbiter_i/n62 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n79  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [4] : \oc8051_xiommu1/oc8051_memarbiter_i/n63 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n80  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [3] : \oc8051_xiommu1/oc8051_memarbiter_i/n64 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n81  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [2] : \oc8051_xiommu1/oc8051_memarbiter_i/n65 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n82  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n66 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n83  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_addr [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n67 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3494 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [15] : \oc8051_xiommu1/oc8051_memarbiter_i/n68 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3478 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [14] : \oc8051_xiommu1/oc8051_memarbiter_i/n69 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3470 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [13] : \oc8051_xiommu1/oc8051_memarbiter_i/n70 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3466 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [12] : \oc8051_xiommu1/oc8051_memarbiter_i/n71 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_1377 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [11] : \oc8051_xiommu1/oc8051_memarbiter_i/n72 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3710 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [10] : \oc8051_xiommu1/oc8051_memarbiter_i/n73 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3706 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [9] : \oc8051_xiommu1/oc8051_memarbiter_i/n74 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_1401 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [8] : \oc8051_xiommu1/oc8051_memarbiter_i/n75 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/addr_out [7] = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [7] : \oc8051_xiommu1/oc8051_memarbiter_i/n76 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/addr_out [6] = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [6] : \oc8051_xiommu1/oc8051_memarbiter_i/n77 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/addr_out [5] = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [5] : \oc8051_xiommu1/oc8051_memarbiter_i/n78 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3986 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [4] : \oc8051_xiommu1/oc8051_memarbiter_i/n79 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3970 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [3] : \oc8051_xiommu1/oc8051_memarbiter_i/n80 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3962 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [2] : \oc8051_xiommu1/oc8051_memarbiter_i/n81 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_3958 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n82 ;   // oc8051_memarbiter.v(139)
    assign _cvpt_1411 = _cvpt_1255 ? \oc8051_xiommu1/proc_addr [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n83 ;   // oc8051_memarbiter.v(139)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n108  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [7] : \oc8051_xiommu1/memwr_xram_data_out [7];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n109  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [6] : \oc8051_xiommu1/memwr_xram_data_out [6];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n110  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [5] : \oc8051_xiommu1/memwr_xram_data_out [5];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n111  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [4] : \oc8051_xiommu1/memwr_xram_data_out [4];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n112  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [3] : \oc8051_xiommu1/memwr_xram_data_out [3];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n113  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [2] : \oc8051_xiommu1/memwr_xram_data_out [2];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n114  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [1] : \oc8051_xiommu1/memwr_xram_data_out [1];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n115  = _cvpt_1252 ? \oc8051_xiommu1/exp_xram_data_out [0] : \oc8051_xiommu1/memwr_xram_data_out [0];   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n116  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [7] : \oc8051_xiommu1/oc8051_memarbiter_i/n108 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n117  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [6] : \oc8051_xiommu1/oc8051_memarbiter_i/n109 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n118  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [5] : \oc8051_xiommu1/oc8051_memarbiter_i/n110 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n119  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [4] : \oc8051_xiommu1/oc8051_memarbiter_i/n111 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n120  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [3] : \oc8051_xiommu1/oc8051_memarbiter_i/n112 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n121  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [2] : \oc8051_xiommu1/oc8051_memarbiter_i/n113 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n122  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n114 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n123  = _cvpt_1253 ? \oc8051_xiommu1/sha_xram_data_out [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n115 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n124  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [7] : \oc8051_xiommu1/oc8051_memarbiter_i/n116 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n125  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [6] : \oc8051_xiommu1/oc8051_memarbiter_i/n117 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n126  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [5] : \oc8051_xiommu1/oc8051_memarbiter_i/n118 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n127  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [4] : \oc8051_xiommu1/oc8051_memarbiter_i/n119 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n128  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [3] : \oc8051_xiommu1/oc8051_memarbiter_i/n120 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n129  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [2] : \oc8051_xiommu1/oc8051_memarbiter_i/n121 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n130  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n122 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n131  = _cvpt_1254 ? \oc8051_xiommu1/aes_xram_data_out [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n123 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [7] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n124 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [6] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n125 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [5] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n126 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [4] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n127 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [3] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n128 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [2] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n129 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [1] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [1] : \oc8051_xiommu1/oc8051_memarbiter_i/n130 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/memarbiter_data_in [0] = _cvpt_1255 ? \oc8051_xiommu1/proc_data_in [0] : \oc8051_xiommu1/oc8051_memarbiter_i/n131 ;   // oc8051_memarbiter.v(144)
    assign \oc8051_xiommu1/proc_ack  = _cvpt_1255 ? \oc8051_xiommu1/ack_in  : 1'b0;   // oc8051_memarbiter.v(146)
    assign _cvpt_392 = _cvpt_1254 ? \oc8051_xiommu1/ack_in  : 1'b0;   // oc8051_memarbiter.v(147)
    assign \oc8051_xiommu1/sha_xram_ack  = _cvpt_1253 ? \oc8051_xiommu1/ack_in  : 1'b0;   // oc8051_memarbiter.v(148)
    assign \oc8051_xiommu1/exp_xram_ack  = _cvpt_1252 ? \oc8051_xiommu1/ack_in  : 1'b0;   // oc8051_memarbiter.v(149)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n152 , \oc8051_xiommu1/selected_port [2]) ;   // oc8051_memarbiter.v(150)
    xor (_cvpt_3401, 1'b0, _cvpt_1411) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/memwr_xram_ack  = _cvpt_1360 ? \oc8051_xiommu1/ack_in  : 1'b0;   // oc8051_memarbiter.v(150)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_inuse_next , \oc8051_xiommu1/ack_in ) ;   // oc8051_memarbiter.v(164)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/n156 , \oc8051_xiommu1/proc_stb , 
        \oc8051_xiommu1/aes_xram_stb ) ;   // oc8051_memarbiter.v(168)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/n157 , \oc8051_xiommu1/oc8051_memarbiter_i/n156 , 
        \oc8051_xiommu1/sha_xram_stb ) ;   // oc8051_memarbiter.v(168)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/n158 , \oc8051_xiommu1/oc8051_memarbiter_i/n157 , 
        \oc8051_xiommu1/exp_xram_stb ) ;   // oc8051_memarbiter.v(168)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/n159 , \oc8051_xiommu1/oc8051_memarbiter_i/n158 , 
        \oc8051_xiommu1/memwr_xram_stb ) ;   // oc8051_memarbiter.v(168)
    and (\oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_idle_next , \oc8051_xiommu1/oc8051_memarbiter_i/n159 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_inuse_next ) ;   // oc8051_memarbiter.v(168)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_next  = _cvpt_1361 ? \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_inuse_next  : \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_idle_next ;   // oc8051_memarbiter.v(172)
    not (_cvpt_1370, _cvpt_1361) ;   // oc8051_memarbiter.v(176)
    and (_cvpt_1367, _cvpt_1370, \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_next ) ;   // oc8051_memarbiter.v(176)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n168 , \oc8051_xiommu1/proc_stb ) ;   // oc8051_memarbiter.v(179)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n169 , \oc8051_xiommu1/aes_xram_stb ) ;   // oc8051_memarbiter.v(179)
    and (\oc8051_xiommu1/oc8051_memarbiter_i/n170 , \oc8051_xiommu1/oc8051_memarbiter_i/n168 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n169 ) ;   // oc8051_memarbiter.v(179)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n171 , \oc8051_xiommu1/sha_xram_stb ) ;   // oc8051_memarbiter.v(179)
    and (\oc8051_xiommu1/oc8051_memarbiter_i/n172 , \oc8051_xiommu1/oc8051_memarbiter_i/n170 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n171 ) ;   // oc8051_memarbiter.v(179)
    not (\oc8051_xiommu1/oc8051_memarbiter_i/n173 , \oc8051_xiommu1/exp_xram_stb ) ;   // oc8051_memarbiter.v(179)
    and (\oc8051_xiommu1/oc8051_memarbiter_i/n174 , \oc8051_xiommu1/oc8051_memarbiter_i/n172 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/n173 ) ;   // oc8051_memarbiter.v(179)
    and (_cvpt_1365, \oc8051_xiommu1/oc8051_memarbiter_i/n174 , \oc8051_xiommu1/memwr_xram_stb ) ;   // oc8051_memarbiter.v(179)
    and (_cvpt_1363, \oc8051_xiommu1/oc8051_memarbiter_i/n172 , \oc8051_xiommu1/exp_xram_stb ) ;   // oc8051_memarbiter.v(180)
    and (_cvpt_1362, \oc8051_xiommu1/oc8051_memarbiter_i/n170 , \oc8051_xiommu1/sha_xram_stb ) ;   // oc8051_memarbiter.v(181)
    and (\oc8051_xiommu1/oc8051_memarbiter_i/n187 , \oc8051_xiommu1/oc8051_memarbiter_i/n168 , 
        \oc8051_xiommu1/aes_xram_stb ) ;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n188  = _cvpt_1362 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/n187 ;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n189  = _cvpt_1363 ? 1'b1 : _cvpt_1362;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n190  = _cvpt_1363 ? 1'b1 : \oc8051_xiommu1/oc8051_memarbiter_i/n188 ;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [1] = _cvpt_1365 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/n189 ;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [0] = _cvpt_1365 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/n190 ;   // oc8051_memarbiter.v(182)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [2] = _cvpt_1367 ? _cvpt_1365 : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [2];   // oc8051_memarbiter.v(185)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [1] = _cvpt_1367 ? \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [1] : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [1];   // oc8051_memarbiter.v(185)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [0] = _cvpt_1367 ? \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [0] : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [0];   // oc8051_memarbiter.v(185)
    assign \oc8051_xiommu1/selected_port [2] = _cvpt_1370 ? _cvpt_1365 : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [2];   // oc8051_memarbiter.v(189)
    assign \oc8051_xiommu1/selected_port [1] = _cvpt_1370 ? \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [1] : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [1];   // oc8051_memarbiter.v(189)
    assign \oc8051_xiommu1/selected_port [0] = _cvpt_1370 ? \oc8051_xiommu1/oc8051_memarbiter_i/arbit_winner [0] : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [0];   // oc8051_memarbiter.v(189)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n201  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/arbiter_state_next ;   // oc8051_memarbiter.v(200)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n202  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [2];   // oc8051_memarbiter.v(200)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n203  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [1];   // oc8051_memarbiter.v(200)
    assign \oc8051_xiommu1/oc8051_memarbiter_i/n204  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder_next [0];   // oc8051_memarbiter.v(200)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_memarbiter_i/i206  (.d(\oc8051_xiommu1/oc8051_memarbiter_i/n202 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [2]));   // oc8051_memarbiter.v(201)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_memarbiter_i/i207  (.d(\oc8051_xiommu1/oc8051_memarbiter_i/n203 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [1]));   // oc8051_memarbiter.v(201)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_memarbiter_i/i208  (.d(\oc8051_xiommu1/oc8051_memarbiter_i/n204 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_memarbiter_i/arbit_holder [0]));   // oc8051_memarbiter.v(201)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_memarbiter_i/i205  (.d(\oc8051_xiommu1/oc8051_memarbiter_i/n201 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(_cvpt_1361));   // oc8051_memarbiter.v(201)
    xor (_cvpt_3417, _cvpt_1411, 1'b1) ;   // oc8051_page_table.v(65)
    xor (_cvpt_3433, 1'b0, _cvpt_1411) ;   // oc8051_page_table.v(66)
    and (_cvpt_1386, \oc8051_xiommu1/oc8051_page_table_i/n4 , \oc8051_xiommu1/oc8051_page_table_i/n5 ) ;   // oc8051_page_table.v(65)
    xor (_cvpt_3449, _cvpt_1411, 1'b1) ;   // oc8051_page_table.v(66)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n1 , _cvpt_1411, 
        _cvpt_3958) ;   // oc8051_page_table.v(70)
    and (_cvpt_1378, \oc8051_xiommu1/oc8051_page_table_i/n7 , \oc8051_xiommu1/oc8051_page_table_i/n8 ) ;   // oc8051_page_table.v(66)
    or (\oc8051_xiommu1/pt_addr_range , _cvpt_1386, _cvpt_1378) ;   // oc8051_page_table.v(67)
    not (\oc8051_xiommu1/oc8051_page_table_i/n11 , \oc8051_xiommu1/addr_out [6]) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n12 , \oc8051_xiommu1/addr_out [7]) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n13 , _cvpt_1401) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n14 , _cvpt_3706) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n15 , _cvpt_3710) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n16 , _cvpt_1377) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n17 , _cvpt_3466) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n18 , _cvpt_3470) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n19 , _cvpt_3478) ;   // oc8051_page_table.v(70)
    not (\oc8051_xiommu1/oc8051_page_table_i/n20 , _cvpt_3494) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n1 , \oc8051_xiommu1/oc8051_page_table_i/n22 , 
        _cvpt_3958) ;   // oc8051_page_table.v(71)
    not (\oc8051_xiommu1/oc8051_page_table_i/n22 , _cvpt_1411) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n1 , _cvpt_1411, 
        \oc8051_xiommu1/oc8051_page_table_i/n34 ) ;   // oc8051_page_table.v(72)
    not (\oc8051_xiommu1/oc8051_page_table_i/n34 , _cvpt_3958) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n1 , \oc8051_xiommu1/oc8051_page_table_i/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/n34 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n1 , _cvpt_1411, 
        _cvpt_3958) ;   // oc8051_page_table.v(74)
    not (\oc8051_xiommu1/oc8051_page_table_i/n59 , _cvpt_3962) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n1 , \oc8051_xiommu1/oc8051_page_table_i/n22 , 
        _cvpt_3958) ;   // oc8051_page_table.v(75)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [7];   // oc8051_page_table.v(87)
    or (\oc8051_xiommu1/oc8051_page_table_i/n84 , _cvpt_3288, _cvpt_3272) ;   // oc8051_page_table.v(76)
    or (\oc8051_xiommu1/oc8051_page_table_i/n85 , \oc8051_xiommu1/oc8051_page_table_i/n84 , 
        _cvpt_3280) ;   // oc8051_page_table.v(76)
    or (\oc8051_xiommu1/oc8051_page_table_i/n86 , \oc8051_xiommu1/oc8051_page_table_i/n85 , 
        _cvpt_3264) ;   // oc8051_page_table.v(76)
    or (\oc8051_xiommu1/oc8051_page_table_i/n87 , \oc8051_xiommu1/oc8051_page_table_i/n86 , 
        \oc8051_xiommu1/oc8051_page_table_i/ia_pc_hi ) ;   // oc8051_page_table.v(76)
    or (\oc8051_xiommu1/ia_addr_range , \oc8051_xiommu1/oc8051_page_table_i/n87 , 
        _cvpt_3256) ;   // oc8051_page_table.v(76)
    and (\oc8051_xiommu1/oc8051_page_table_i/n89 , \oc8051_xiommu1/priv_lvl , 
        _cvpt_119) ;   // oc8051_page_table.v(79)
    and (_cvpt_1420, \oc8051_xiommu1/oc8051_page_table_i/n89 , _cvpt_1386) ;   // oc8051_page_table.v(79)
    and (_cvpt_1435, \oc8051_xiommu1/oc8051_page_table_i/n89 , _cvpt_1378) ;   // oc8051_page_table.v(80)
    assign \oc8051_xiommu1/oc8051_page_table_i/n93  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [7] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n94  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [6] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n95  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [5] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n96  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [4] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n97  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [3] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n98  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [2] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n99  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [1] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/n100  = _cvpt_1378 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [0] : 1'b0;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [7] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [7] : \oc8051_xiommu1/oc8051_page_table_i/n93 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [6] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [6] : \oc8051_xiommu1/oc8051_page_table_i/n94 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [5] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [5] : \oc8051_xiommu1/oc8051_page_table_i/n95 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [4] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [4] : \oc8051_xiommu1/oc8051_page_table_i/n96 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [3] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [3] : \oc8051_xiommu1/oc8051_page_table_i/n97 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [2] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [2] : \oc8051_xiommu1/oc8051_page_table_i/n98 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [1] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [1] : \oc8051_xiommu1/oc8051_page_table_i/n99 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/data_out_pt [0] = _cvpt_1386 ? \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [0] : \oc8051_xiommu1/oc8051_page_table_i/n100 ;   // oc8051_page_table.v(84)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n1  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n115  : \oc8051_xiommu1/oc8051_page_table_i/n116 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n1  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n1  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n124  : \oc8051_xiommu1/oc8051_page_table_i/n125 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [7];   // oc8051_page_table.v(92)
    and (\oc8051_xiommu1/ack_pt , _cvpt_119, \oc8051_xiommu1/pt_addr_range ) ;   // oc8051_page_table.v(89)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [7] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n128  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [6] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n129  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [5] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n130  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [4] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n131  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [3] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n132  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [2] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n133  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [1] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n134  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_wr [0] = _cvpt_1420 ? \oc8051_xiommu1/oc8051_page_table_i/n135  : 1'b0;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n1  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0];   // oc8051_page_table.v(93)
    not (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n8 , _cvpt_1411) ;   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [7] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n144  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [6] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n145  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [5] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n146  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [4] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n147  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [3] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n148  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [2] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n149  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [1] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n150  : 1'b0;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/data_out_rd [0] = _cvpt_1435 ? \oc8051_xiommu1/oc8051_page_table_i/n151  : 1'b0;   // oc8051_page_table.v(93)
    and (_cvpt_2211, \oc8051_xiommu1/write_pt , _cvpt_1420) ;   // oc8051_page_table.v(106)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_or_2475/n1 , \oc8051_xiommu1/selected_port [1], 
        \oc8051_xiommu1/selected_port [2]) ;   // oc8051_page_table.v(129)
    assign \oc8051_xiommu1/oc8051_page_table_i/n194  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n195  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n196  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n197  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n198  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n199  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n200  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n201  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n202  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n203  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n204  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n205  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n206  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n207  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n208  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n209  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n210  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n211  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n212  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n213  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n214  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n215  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n216  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n217  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n218  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n219  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n220  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n221  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n222  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n223  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n224  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n225  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n226  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n227  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n228  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n229  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n230  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n231  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n232  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n233  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n234  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n235  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n236  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n237  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n238  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n239  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n240  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n241  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n242  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n243  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n244  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n245  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n246  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n247  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n248  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n249  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n250  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n251  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n252  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n253  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n254  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n255  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n256  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n257  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n258  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n259  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n260  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n261  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n262  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n263  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n264  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n265  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n266  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n267  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n268  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n269  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n270  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n271  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n272  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n273  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n274  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n275  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n276  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n277  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n278  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n279  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n280  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n281  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n282  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n283  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n284  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n285  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n286  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n287  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n288  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n289  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n290  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n291  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n292  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n293  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n294  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n295  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n296  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n297  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n298  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n299  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n300  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n301  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n302  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n303  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n304  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n305  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n306  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n307  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n308  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n309  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n310  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n311  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n312  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n313  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n314  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n315  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n316  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n317  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n318  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n319  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n320  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n321  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n322  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n323  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n324  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n325  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n326  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n327  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n328  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n329  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n330  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n331  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n332  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n333  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n334  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n335  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n336  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n337  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n338  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n339  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n340  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n341  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n342  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n343  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n344  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n345  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n346  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n347  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n348  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n349  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n350  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n351  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n352  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n353  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n354  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n355  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n356  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n357  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n358  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n359  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n360  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n361  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n362  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n363  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n364  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n365  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n366  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n367  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n368  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n369  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n370  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n371  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n372  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n373  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n374  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n375  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n376  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n377  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n378  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n379  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n380  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n381  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n382  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n383  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n384  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n385  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n386  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n387  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n388  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n389  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n390  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n391  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n392  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n393  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n394  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n395  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n396  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n397  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n398  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n399  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n400  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n401  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n402  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n403  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n404  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n405  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n406  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n407  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n408  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n409  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n410  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n411  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n412  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n413  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n414  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n415  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n416  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n417  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n418  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n419  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n420  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n421  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n422  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n423  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n424  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n425  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n426  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n427  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n428  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n429  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n430  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n431  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n432  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n433  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n434  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n435  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n436  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n437  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n438  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n439  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n440  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n441  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [0];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n442  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [7];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n443  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [6];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n444  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [5];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n445  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [4];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n446  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [3];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n447  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [2];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n448  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [1];   // oc8051_page_table.v(107)
    assign \oc8051_xiommu1/oc8051_page_table_i/n449  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [0];   // oc8051_page_table.v(107)
    and (_cvpt_1955, \oc8051_xiommu1/write_pt , _cvpt_1435) ;   // oc8051_page_table.v(109)
    assign \oc8051_xiommu1/oc8051_page_table_i/n483  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n484  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n485  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n486  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n487  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n488  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n489  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n490  = _cvpt_1443 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n491  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n492  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n493  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n494  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n495  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n496  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n497  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n498  = _cvpt_1451 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n499  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n500  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n501  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n502  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n503  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n504  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n505  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n506  = _cvpt_1459 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n507  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n508  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n509  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n510  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n511  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n512  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n513  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n514  = _cvpt_1467 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n515  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n516  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n517  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n518  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n519  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n520  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n521  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n522  = _cvpt_1475 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n523  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n524  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n525  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n526  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n527  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n528  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n529  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n530  = _cvpt_1483 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n531  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n532  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n533  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n534  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n535  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n536  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n537  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n538  = _cvpt_1491 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n539  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n540  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n541  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n542  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n543  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n544  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n545  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n546  = _cvpt_1499 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n547  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n548  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n549  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n550  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n551  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n552  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n553  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n554  = _cvpt_1507 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n555  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n556  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n557  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n558  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n559  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n560  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n561  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n562  = _cvpt_1515 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n563  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n564  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n565  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n566  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n567  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n568  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n569  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n570  = _cvpt_1523 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n571  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n572  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n573  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n574  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n575  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n576  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n577  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n578  = _cvpt_1531 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n579  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n580  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n581  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n582  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n583  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n584  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n585  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n586  = _cvpt_1539 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n587  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n588  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n589  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n590  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n591  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n592  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n593  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n594  = _cvpt_1547 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n595  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n596  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n597  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n598  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n599  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n600  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n601  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n602  = _cvpt_1555 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n603  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n604  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n605  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n606  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n607  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n608  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n609  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n610  = _cvpt_1563 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n611  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n612  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n613  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n614  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n615  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n616  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n617  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n618  = _cvpt_1571 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n619  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n620  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n621  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n622  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n623  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n624  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n625  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n626  = _cvpt_1579 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n627  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n628  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n629  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n630  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n631  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n632  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n633  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n634  = _cvpt_1587 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n635  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n636  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n637  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n638  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n639  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n640  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n641  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n642  = _cvpt_1595 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n643  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n644  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n645  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n646  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n647  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n648  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n649  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n650  = _cvpt_1603 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n651  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n652  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n653  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n654  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n655  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n656  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n657  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n658  = _cvpt_1611 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n659  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n660  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n661  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n662  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n663  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n664  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n665  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n666  = _cvpt_1619 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n667  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n668  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n669  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n670  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n671  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n672  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n673  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n674  = _cvpt_1627 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n675  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n676  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n677  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n678  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n679  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n680  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n681  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n682  = _cvpt_1635 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n683  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n684  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n685  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n686  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n687  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n688  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n689  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n690  = _cvpt_1643 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n691  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n692  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n693  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n694  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n695  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n696  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n697  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n698  = _cvpt_1651 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n699  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n700  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n701  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n702  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n703  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n704  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n705  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n706  = _cvpt_1659 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n707  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n708  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n709  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n710  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n711  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n712  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n713  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n714  = _cvpt_1667 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n715  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n716  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n717  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n718  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n719  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n720  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n721  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n722  = _cvpt_1675 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n723  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n724  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n725  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n726  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n727  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n728  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n729  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n730  = _cvpt_1683 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n731  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n732  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n733  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n734  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n735  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n736  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n737  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n738  = _cvpt_1691 ? \oc8051_xiommu1/memarbiter_data_in [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0];   // oc8051_page_table.v(110)
    assign \oc8051_xiommu1/oc8051_page_table_i/n739  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n483  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n740  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n484  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n741  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n485  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n742  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n486  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n743  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n487  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n744  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n488  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n745  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n489  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n746  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n490  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n747  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n491  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n748  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n492  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n749  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n493  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n750  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n494  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n751  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n495  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n752  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n496  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n753  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n497  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n754  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n498  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n755  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n499  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n756  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n500  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n757  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n501  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n758  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n502  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n759  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n503  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n760  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n504  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n761  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n505  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n762  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n506  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n763  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n507  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n764  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n508  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n765  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n509  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n766  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n510  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n767  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n511  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n768  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n512  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n769  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n513  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n770  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n514  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n771  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n515  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n772  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n516  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n773  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n517  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n774  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n518  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n775  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n519  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n776  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n520  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n777  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n521  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n778  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n522  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n779  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n523  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n780  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n524  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n781  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n525  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n782  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n526  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n783  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n527  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n784  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n528  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n785  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n529  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n786  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n530  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n787  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n531  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n788  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n532  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n789  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n533  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n790  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n534  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n791  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n535  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n792  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n536  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n793  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n537  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n794  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n538  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n795  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n539  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n796  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n540  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n797  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n541  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n798  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n542  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n799  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n543  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n800  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n544  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n801  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n545  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n802  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n546  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n803  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n547  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n804  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n548  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n805  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n549  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n806  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n550  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n807  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n551  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n808  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n552  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n809  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n553  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n810  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n554  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n811  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n555  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n812  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n556  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n813  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n557  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n814  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n558  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n815  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n559  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n816  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n560  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n817  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n561  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n818  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n562  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n819  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n563  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n820  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n564  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n821  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n565  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n822  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n566  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n823  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n567  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n824  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n568  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n825  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n569  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n826  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n570  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n827  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n571  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n828  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n572  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n829  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n573  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n830  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n574  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n831  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n575  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n832  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n576  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n833  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n577  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n834  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n578  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n835  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n579  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n836  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n580  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n837  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n581  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n838  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n582  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n839  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n583  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n840  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n584  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n841  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n585  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n842  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n586  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n843  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n587  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n844  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n588  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n845  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n589  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n846  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n590  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n847  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n591  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n848  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n592  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n849  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n593  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n850  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n594  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n851  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n595  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n852  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n596  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n853  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n597  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n854  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n598  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n855  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n599  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n856  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n600  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n857  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n601  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n858  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n602  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n859  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n603  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n860  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n604  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n861  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n605  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n862  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n606  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n863  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n607  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n864  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n608  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n865  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n609  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n866  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n610  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n867  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n611  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n868  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n612  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n869  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n613  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n870  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n614  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n871  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n615  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n872  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n616  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n873  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n617  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n874  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n618  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n875  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n619  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n876  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n620  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n877  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n621  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n878  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n622  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n879  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n623  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n880  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n624  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n881  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n625  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n882  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n626  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n883  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n627  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n884  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n628  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n885  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n629  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n886  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n630  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n887  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n631  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n888  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n632  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n889  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n633  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n890  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n634  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n891  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n635  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n892  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n636  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n893  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n637  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n894  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n638  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n895  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n639  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n896  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n640  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n897  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n641  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n898  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n642  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n899  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n643  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n900  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n644  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n901  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n645  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n902  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n646  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n903  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n647  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n904  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n648  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n905  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n649  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n906  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n650  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n907  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n651  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n908  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n652  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n909  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n653  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n910  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n654  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n911  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n655  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n912  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n656  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n913  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n657  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n914  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n658  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n915  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n659  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n916  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n660  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n917  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n661  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n918  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n662  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n919  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n663  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n920  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n664  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n921  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n665  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n922  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n666  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n923  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n667  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n924  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n668  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n925  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n669  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n926  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n670  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n927  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n671  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n928  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n672  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n929  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n673  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n930  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n674  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n931  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n675  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n932  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n676  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n933  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n677  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n934  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n678  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n935  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n679  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n936  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n680  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n937  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n681  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n938  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n682  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n939  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n683  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n940  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n684  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n941  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n685  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n942  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n686  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n943  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n687  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n944  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n688  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n945  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n689  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n946  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n690  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n947  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n691  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n948  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n692  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n949  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n693  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n950  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n694  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n951  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n695  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n952  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n696  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n953  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n697  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n954  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n698  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n955  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n699  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n956  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n700  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n957  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n701  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n958  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n702  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n959  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n703  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n960  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n704  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n961  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n705  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n962  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n706  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n963  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n707  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n964  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n708  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n965  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n709  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n966  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n710  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n967  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n711  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n968  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n712  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n969  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n713  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n970  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n714  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n971  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n715  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n972  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n716  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n973  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n717  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n974  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n718  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n975  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n719  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n976  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n720  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n977  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n721  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n978  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n722  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n979  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n723  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n980  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n724  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n981  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n725  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n982  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n726  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n983  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n727  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n984  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n728  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n985  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n729  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n986  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n730  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n987  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n731  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n988  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n732  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n989  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n733  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n990  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n734  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n991  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n735  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n992  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n736  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n993  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n737  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n994  = _cvpt_1955 ? \oc8051_xiommu1/oc8051_page_table_i/n738  : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n995  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n194  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n996  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n195  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n997  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n196  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n998  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n197  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n999  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n198  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1000  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n199  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1001  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n200  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1002  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n201  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1003  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n202  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1004  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n203  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1005  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n204  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1006  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n205  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1007  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n206  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1008  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n207  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1009  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n208  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1010  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n209  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1011  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n210  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1012  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n211  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1013  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n212  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1014  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n213  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1015  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n214  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1016  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n215  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1017  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n216  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1018  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n217  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1019  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n218  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1020  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n219  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1021  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n220  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1022  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n221  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1023  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n222  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1024  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n223  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1025  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n224  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1026  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n225  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1027  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n226  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1028  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n227  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1029  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n228  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1030  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n229  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1031  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n230  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1032  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n231  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1033  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n232  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1034  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n233  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1035  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n234  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1036  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n235  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1037  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n236  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1038  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n237  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1039  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n238  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1040  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n239  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1041  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n240  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1042  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n241  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1043  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n242  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1044  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n243  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1045  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n244  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1046  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n245  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1047  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n246  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1048  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n247  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1049  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n248  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1050  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n249  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1051  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n250  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1052  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n251  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1053  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n252  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1054  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n253  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1055  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n254  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1056  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n255  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1057  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n256  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1058  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n257  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1059  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n258  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1060  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n259  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1061  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n260  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1062  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n261  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1063  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n262  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1064  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n263  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1065  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n264  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1066  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n265  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1067  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n266  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1068  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n267  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1069  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n268  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1070  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n269  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1071  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n270  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1072  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n271  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1073  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n272  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1074  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n273  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1075  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n274  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1076  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n275  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1077  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n276  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1078  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n277  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1079  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n278  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1080  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n279  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1081  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n280  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1082  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n281  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1083  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n282  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1084  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n283  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1085  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n284  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1086  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n285  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1087  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n286  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1088  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n287  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1089  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n288  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1090  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n289  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1091  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n290  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1092  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n291  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1093  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n292  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1094  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n293  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1095  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n294  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1096  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n295  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1097  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n296  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1098  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n297  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1099  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n298  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1100  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n299  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1101  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n300  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1102  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n301  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1103  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n302  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1104  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n303  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1105  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n304  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1106  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n305  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1107  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n306  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1108  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n307  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1109  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n308  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1110  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n309  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1111  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n310  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1112  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n311  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1113  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n312  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1114  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n313  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1115  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n314  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1116  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n315  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1117  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n316  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1118  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n317  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1119  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n318  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1120  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n319  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1121  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n320  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1122  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n321  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1123  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n322  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1124  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n323  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1125  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n324  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1126  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n325  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1127  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n326  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1128  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n327  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1129  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n328  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1130  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n329  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1131  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n330  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1132  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n331  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1133  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n332  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1134  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n333  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1135  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n334  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1136  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n335  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1137  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n336  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1138  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n337  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1139  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n338  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1140  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n339  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1141  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n340  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1142  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n341  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1143  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n342  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1144  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n343  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1145  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n344  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1146  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n345  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1147  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n346  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1148  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n347  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1149  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n348  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1150  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n349  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1151  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n350  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1152  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n351  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1153  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n352  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1154  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n353  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1155  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n354  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1156  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n355  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1157  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n356  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1158  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n357  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1159  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n358  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1160  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n359  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1161  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n360  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1162  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n361  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1163  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n362  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1164  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n363  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1165  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n364  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1166  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n365  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1167  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n366  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1168  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n367  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1169  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n368  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1170  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n369  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1171  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n370  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1172  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n371  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1173  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n372  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1174  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n373  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1175  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n374  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1176  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n375  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1177  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n376  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1178  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n377  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1179  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n378  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1180  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n379  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1181  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n380  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1182  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n381  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1183  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n382  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1184  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n383  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1185  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n384  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1186  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n385  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1187  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n386  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1188  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n387  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1189  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n388  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1190  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n389  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1191  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n390  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1192  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n391  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1193  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n392  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1194  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n393  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1195  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n394  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1196  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n395  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1197  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n396  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1198  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n397  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1199  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n398  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1200  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n399  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1201  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n400  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1202  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n401  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1203  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n402  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1204  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n403  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1205  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n404  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1206  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n405  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1207  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n406  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1208  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n407  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1209  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n408  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1210  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n409  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1211  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n410  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1212  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n411  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1213  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n412  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1214  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n413  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1215  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n414  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1216  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n415  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1217  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n416  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1218  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n417  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1219  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n418  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1220  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n419  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1221  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n420  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1222  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n421  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1223  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n422  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1224  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n423  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1225  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n424  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1226  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n425  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1227  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n426  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1228  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n427  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1229  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n428  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1230  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n429  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1231  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n430  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1232  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n431  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1233  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n432  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1234  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n433  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1235  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n434  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1236  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n435  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1237  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n436  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1238  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n437  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1239  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n438  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1240  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n439  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1241  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n440  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1242  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n441  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1243  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n442  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [7];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1244  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n443  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [6];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1245  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n444  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [5];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1246  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n445  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [4];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1247  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n446  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [3];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1248  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n447  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [2];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1249  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n448  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [1];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1250  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/n449  : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [0];   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1251  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7] : \oc8051_xiommu1/oc8051_page_table_i/n739 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1252  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6] : \oc8051_xiommu1/oc8051_page_table_i/n740 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1253  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5] : \oc8051_xiommu1/oc8051_page_table_i/n741 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1254  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4] : \oc8051_xiommu1/oc8051_page_table_i/n742 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1255  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3] : \oc8051_xiommu1/oc8051_page_table_i/n743 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1256  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2] : \oc8051_xiommu1/oc8051_page_table_i/n744 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1257  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1] : \oc8051_xiommu1/oc8051_page_table_i/n745 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1258  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0] : \oc8051_xiommu1/oc8051_page_table_i/n746 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1259  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7] : \oc8051_xiommu1/oc8051_page_table_i/n747 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1260  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6] : \oc8051_xiommu1/oc8051_page_table_i/n748 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1261  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5] : \oc8051_xiommu1/oc8051_page_table_i/n749 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1262  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4] : \oc8051_xiommu1/oc8051_page_table_i/n750 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1263  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3] : \oc8051_xiommu1/oc8051_page_table_i/n751 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1264  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2] : \oc8051_xiommu1/oc8051_page_table_i/n752 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1265  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1] : \oc8051_xiommu1/oc8051_page_table_i/n753 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1266  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0] : \oc8051_xiommu1/oc8051_page_table_i/n754 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1267  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7] : \oc8051_xiommu1/oc8051_page_table_i/n755 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1268  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6] : \oc8051_xiommu1/oc8051_page_table_i/n756 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1269  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5] : \oc8051_xiommu1/oc8051_page_table_i/n757 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1270  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4] : \oc8051_xiommu1/oc8051_page_table_i/n758 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1271  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3] : \oc8051_xiommu1/oc8051_page_table_i/n759 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1272  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2] : \oc8051_xiommu1/oc8051_page_table_i/n760 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1273  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1] : \oc8051_xiommu1/oc8051_page_table_i/n761 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1274  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0] : \oc8051_xiommu1/oc8051_page_table_i/n762 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1275  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7] : \oc8051_xiommu1/oc8051_page_table_i/n763 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1276  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6] : \oc8051_xiommu1/oc8051_page_table_i/n764 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1277  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5] : \oc8051_xiommu1/oc8051_page_table_i/n765 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1278  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4] : \oc8051_xiommu1/oc8051_page_table_i/n766 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1279  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3] : \oc8051_xiommu1/oc8051_page_table_i/n767 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1280  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2] : \oc8051_xiommu1/oc8051_page_table_i/n768 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1281  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1] : \oc8051_xiommu1/oc8051_page_table_i/n769 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1282  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0] : \oc8051_xiommu1/oc8051_page_table_i/n770 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1283  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7] : \oc8051_xiommu1/oc8051_page_table_i/n771 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1284  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6] : \oc8051_xiommu1/oc8051_page_table_i/n772 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1285  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5] : \oc8051_xiommu1/oc8051_page_table_i/n773 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1286  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4] : \oc8051_xiommu1/oc8051_page_table_i/n774 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1287  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3] : \oc8051_xiommu1/oc8051_page_table_i/n775 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1288  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2] : \oc8051_xiommu1/oc8051_page_table_i/n776 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1289  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1] : \oc8051_xiommu1/oc8051_page_table_i/n777 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1290  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0] : \oc8051_xiommu1/oc8051_page_table_i/n778 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1291  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7] : \oc8051_xiommu1/oc8051_page_table_i/n779 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1292  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6] : \oc8051_xiommu1/oc8051_page_table_i/n780 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1293  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5] : \oc8051_xiommu1/oc8051_page_table_i/n781 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1294  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4] : \oc8051_xiommu1/oc8051_page_table_i/n782 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1295  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3] : \oc8051_xiommu1/oc8051_page_table_i/n783 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1296  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2] : \oc8051_xiommu1/oc8051_page_table_i/n784 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1297  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1] : \oc8051_xiommu1/oc8051_page_table_i/n785 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1298  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0] : \oc8051_xiommu1/oc8051_page_table_i/n786 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1299  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7] : \oc8051_xiommu1/oc8051_page_table_i/n787 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1300  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6] : \oc8051_xiommu1/oc8051_page_table_i/n788 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1301  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5] : \oc8051_xiommu1/oc8051_page_table_i/n789 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1302  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4] : \oc8051_xiommu1/oc8051_page_table_i/n790 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1303  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3] : \oc8051_xiommu1/oc8051_page_table_i/n791 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1304  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2] : \oc8051_xiommu1/oc8051_page_table_i/n792 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1305  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1] : \oc8051_xiommu1/oc8051_page_table_i/n793 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1306  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0] : \oc8051_xiommu1/oc8051_page_table_i/n794 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1307  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7] : \oc8051_xiommu1/oc8051_page_table_i/n795 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1308  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6] : \oc8051_xiommu1/oc8051_page_table_i/n796 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1309  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5] : \oc8051_xiommu1/oc8051_page_table_i/n797 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1310  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4] : \oc8051_xiommu1/oc8051_page_table_i/n798 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1311  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3] : \oc8051_xiommu1/oc8051_page_table_i/n799 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1312  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2] : \oc8051_xiommu1/oc8051_page_table_i/n800 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1313  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1] : \oc8051_xiommu1/oc8051_page_table_i/n801 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1314  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0] : \oc8051_xiommu1/oc8051_page_table_i/n802 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1315  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7] : \oc8051_xiommu1/oc8051_page_table_i/n803 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1316  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6] : \oc8051_xiommu1/oc8051_page_table_i/n804 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1317  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5] : \oc8051_xiommu1/oc8051_page_table_i/n805 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1318  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4] : \oc8051_xiommu1/oc8051_page_table_i/n806 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1319  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3] : \oc8051_xiommu1/oc8051_page_table_i/n807 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1320  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2] : \oc8051_xiommu1/oc8051_page_table_i/n808 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1321  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1] : \oc8051_xiommu1/oc8051_page_table_i/n809 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1322  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0] : \oc8051_xiommu1/oc8051_page_table_i/n810 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1323  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7] : \oc8051_xiommu1/oc8051_page_table_i/n811 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1324  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6] : \oc8051_xiommu1/oc8051_page_table_i/n812 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1325  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5] : \oc8051_xiommu1/oc8051_page_table_i/n813 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1326  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4] : \oc8051_xiommu1/oc8051_page_table_i/n814 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1327  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3] : \oc8051_xiommu1/oc8051_page_table_i/n815 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1328  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2] : \oc8051_xiommu1/oc8051_page_table_i/n816 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1329  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1] : \oc8051_xiommu1/oc8051_page_table_i/n817 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1330  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0] : \oc8051_xiommu1/oc8051_page_table_i/n818 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1331  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7] : \oc8051_xiommu1/oc8051_page_table_i/n819 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1332  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6] : \oc8051_xiommu1/oc8051_page_table_i/n820 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1333  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5] : \oc8051_xiommu1/oc8051_page_table_i/n821 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1334  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4] : \oc8051_xiommu1/oc8051_page_table_i/n822 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1335  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3] : \oc8051_xiommu1/oc8051_page_table_i/n823 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1336  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2] : \oc8051_xiommu1/oc8051_page_table_i/n824 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1337  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1] : \oc8051_xiommu1/oc8051_page_table_i/n825 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1338  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0] : \oc8051_xiommu1/oc8051_page_table_i/n826 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1339  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7] : \oc8051_xiommu1/oc8051_page_table_i/n827 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1340  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6] : \oc8051_xiommu1/oc8051_page_table_i/n828 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1341  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5] : \oc8051_xiommu1/oc8051_page_table_i/n829 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1342  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4] : \oc8051_xiommu1/oc8051_page_table_i/n830 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1343  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3] : \oc8051_xiommu1/oc8051_page_table_i/n831 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1344  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2] : \oc8051_xiommu1/oc8051_page_table_i/n832 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1345  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1] : \oc8051_xiommu1/oc8051_page_table_i/n833 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1346  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0] : \oc8051_xiommu1/oc8051_page_table_i/n834 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1347  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7] : \oc8051_xiommu1/oc8051_page_table_i/n835 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1348  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6] : \oc8051_xiommu1/oc8051_page_table_i/n836 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1349  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5] : \oc8051_xiommu1/oc8051_page_table_i/n837 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1350  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4] : \oc8051_xiommu1/oc8051_page_table_i/n838 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1351  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3] : \oc8051_xiommu1/oc8051_page_table_i/n839 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1352  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2] : \oc8051_xiommu1/oc8051_page_table_i/n840 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1353  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1] : \oc8051_xiommu1/oc8051_page_table_i/n841 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1354  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0] : \oc8051_xiommu1/oc8051_page_table_i/n842 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1355  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7] : \oc8051_xiommu1/oc8051_page_table_i/n843 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1356  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6] : \oc8051_xiommu1/oc8051_page_table_i/n844 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1357  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5] : \oc8051_xiommu1/oc8051_page_table_i/n845 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1358  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4] : \oc8051_xiommu1/oc8051_page_table_i/n846 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1359  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3] : \oc8051_xiommu1/oc8051_page_table_i/n847 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1360  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2] : \oc8051_xiommu1/oc8051_page_table_i/n848 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1361  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1] : \oc8051_xiommu1/oc8051_page_table_i/n849 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1362  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0] : \oc8051_xiommu1/oc8051_page_table_i/n850 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1363  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7] : \oc8051_xiommu1/oc8051_page_table_i/n851 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1364  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6] : \oc8051_xiommu1/oc8051_page_table_i/n852 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1365  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5] : \oc8051_xiommu1/oc8051_page_table_i/n853 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1366  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4] : \oc8051_xiommu1/oc8051_page_table_i/n854 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1367  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3] : \oc8051_xiommu1/oc8051_page_table_i/n855 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1368  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2] : \oc8051_xiommu1/oc8051_page_table_i/n856 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1369  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1] : \oc8051_xiommu1/oc8051_page_table_i/n857 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1370  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0] : \oc8051_xiommu1/oc8051_page_table_i/n858 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1371  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7] : \oc8051_xiommu1/oc8051_page_table_i/n859 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1372  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6] : \oc8051_xiommu1/oc8051_page_table_i/n860 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1373  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5] : \oc8051_xiommu1/oc8051_page_table_i/n861 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1374  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4] : \oc8051_xiommu1/oc8051_page_table_i/n862 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1375  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3] : \oc8051_xiommu1/oc8051_page_table_i/n863 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1376  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2] : \oc8051_xiommu1/oc8051_page_table_i/n864 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1377  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1] : \oc8051_xiommu1/oc8051_page_table_i/n865 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1378  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0] : \oc8051_xiommu1/oc8051_page_table_i/n866 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1379  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7] : \oc8051_xiommu1/oc8051_page_table_i/n867 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1380  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6] : \oc8051_xiommu1/oc8051_page_table_i/n868 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1381  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5] : \oc8051_xiommu1/oc8051_page_table_i/n869 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1382  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4] : \oc8051_xiommu1/oc8051_page_table_i/n870 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1383  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3] : \oc8051_xiommu1/oc8051_page_table_i/n871 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1384  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2] : \oc8051_xiommu1/oc8051_page_table_i/n872 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1385  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1] : \oc8051_xiommu1/oc8051_page_table_i/n873 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1386  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0] : \oc8051_xiommu1/oc8051_page_table_i/n874 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1387  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7] : \oc8051_xiommu1/oc8051_page_table_i/n875 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1388  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6] : \oc8051_xiommu1/oc8051_page_table_i/n876 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1389  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5] : \oc8051_xiommu1/oc8051_page_table_i/n877 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1390  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4] : \oc8051_xiommu1/oc8051_page_table_i/n878 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1391  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3] : \oc8051_xiommu1/oc8051_page_table_i/n879 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1392  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2] : \oc8051_xiommu1/oc8051_page_table_i/n880 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1393  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1] : \oc8051_xiommu1/oc8051_page_table_i/n881 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1394  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0] : \oc8051_xiommu1/oc8051_page_table_i/n882 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1395  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7] : \oc8051_xiommu1/oc8051_page_table_i/n883 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1396  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6] : \oc8051_xiommu1/oc8051_page_table_i/n884 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1397  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5] : \oc8051_xiommu1/oc8051_page_table_i/n885 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1398  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4] : \oc8051_xiommu1/oc8051_page_table_i/n886 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1399  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3] : \oc8051_xiommu1/oc8051_page_table_i/n887 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1400  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2] : \oc8051_xiommu1/oc8051_page_table_i/n888 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1401  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1] : \oc8051_xiommu1/oc8051_page_table_i/n889 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1402  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0] : \oc8051_xiommu1/oc8051_page_table_i/n890 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1403  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7] : \oc8051_xiommu1/oc8051_page_table_i/n891 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1404  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6] : \oc8051_xiommu1/oc8051_page_table_i/n892 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1405  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5] : \oc8051_xiommu1/oc8051_page_table_i/n893 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1406  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4] : \oc8051_xiommu1/oc8051_page_table_i/n894 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1407  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3] : \oc8051_xiommu1/oc8051_page_table_i/n895 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1408  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2] : \oc8051_xiommu1/oc8051_page_table_i/n896 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1409  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1] : \oc8051_xiommu1/oc8051_page_table_i/n897 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1410  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0] : \oc8051_xiommu1/oc8051_page_table_i/n898 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1411  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7] : \oc8051_xiommu1/oc8051_page_table_i/n899 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1412  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6] : \oc8051_xiommu1/oc8051_page_table_i/n900 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1413  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5] : \oc8051_xiommu1/oc8051_page_table_i/n901 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1414  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4] : \oc8051_xiommu1/oc8051_page_table_i/n902 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1415  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3] : \oc8051_xiommu1/oc8051_page_table_i/n903 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1416  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2] : \oc8051_xiommu1/oc8051_page_table_i/n904 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1417  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1] : \oc8051_xiommu1/oc8051_page_table_i/n905 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1418  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0] : \oc8051_xiommu1/oc8051_page_table_i/n906 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1419  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7] : \oc8051_xiommu1/oc8051_page_table_i/n907 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1420  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6] : \oc8051_xiommu1/oc8051_page_table_i/n908 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1421  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5] : \oc8051_xiommu1/oc8051_page_table_i/n909 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1422  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4] : \oc8051_xiommu1/oc8051_page_table_i/n910 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1423  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3] : \oc8051_xiommu1/oc8051_page_table_i/n911 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1424  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2] : \oc8051_xiommu1/oc8051_page_table_i/n912 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1425  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1] : \oc8051_xiommu1/oc8051_page_table_i/n913 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1426  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0] : \oc8051_xiommu1/oc8051_page_table_i/n914 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1427  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7] : \oc8051_xiommu1/oc8051_page_table_i/n915 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1428  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6] : \oc8051_xiommu1/oc8051_page_table_i/n916 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1429  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5] : \oc8051_xiommu1/oc8051_page_table_i/n917 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1430  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4] : \oc8051_xiommu1/oc8051_page_table_i/n918 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1431  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3] : \oc8051_xiommu1/oc8051_page_table_i/n919 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1432  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2] : \oc8051_xiommu1/oc8051_page_table_i/n920 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1433  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1] : \oc8051_xiommu1/oc8051_page_table_i/n921 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1434  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0] : \oc8051_xiommu1/oc8051_page_table_i/n922 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1435  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7] : \oc8051_xiommu1/oc8051_page_table_i/n923 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1436  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6] : \oc8051_xiommu1/oc8051_page_table_i/n924 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1437  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5] : \oc8051_xiommu1/oc8051_page_table_i/n925 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1438  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4] : \oc8051_xiommu1/oc8051_page_table_i/n926 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1439  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3] : \oc8051_xiommu1/oc8051_page_table_i/n927 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1440  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2] : \oc8051_xiommu1/oc8051_page_table_i/n928 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1441  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1] : \oc8051_xiommu1/oc8051_page_table_i/n929 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1442  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0] : \oc8051_xiommu1/oc8051_page_table_i/n930 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1443  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7] : \oc8051_xiommu1/oc8051_page_table_i/n931 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1444  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6] : \oc8051_xiommu1/oc8051_page_table_i/n932 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1445  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5] : \oc8051_xiommu1/oc8051_page_table_i/n933 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1446  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4] : \oc8051_xiommu1/oc8051_page_table_i/n934 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1447  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3] : \oc8051_xiommu1/oc8051_page_table_i/n935 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1448  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2] : \oc8051_xiommu1/oc8051_page_table_i/n936 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1449  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1] : \oc8051_xiommu1/oc8051_page_table_i/n937 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1450  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0] : \oc8051_xiommu1/oc8051_page_table_i/n938 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1451  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7] : \oc8051_xiommu1/oc8051_page_table_i/n939 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1452  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6] : \oc8051_xiommu1/oc8051_page_table_i/n940 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1453  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5] : \oc8051_xiommu1/oc8051_page_table_i/n941 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1454  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4] : \oc8051_xiommu1/oc8051_page_table_i/n942 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1455  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3] : \oc8051_xiommu1/oc8051_page_table_i/n943 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1456  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2] : \oc8051_xiommu1/oc8051_page_table_i/n944 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1457  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1] : \oc8051_xiommu1/oc8051_page_table_i/n945 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1458  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0] : \oc8051_xiommu1/oc8051_page_table_i/n946 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1459  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7] : \oc8051_xiommu1/oc8051_page_table_i/n947 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1460  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6] : \oc8051_xiommu1/oc8051_page_table_i/n948 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1461  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5] : \oc8051_xiommu1/oc8051_page_table_i/n949 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1462  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4] : \oc8051_xiommu1/oc8051_page_table_i/n950 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1463  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3] : \oc8051_xiommu1/oc8051_page_table_i/n951 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1464  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2] : \oc8051_xiommu1/oc8051_page_table_i/n952 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1465  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1] : \oc8051_xiommu1/oc8051_page_table_i/n953 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1466  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0] : \oc8051_xiommu1/oc8051_page_table_i/n954 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1467  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7] : \oc8051_xiommu1/oc8051_page_table_i/n955 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1468  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6] : \oc8051_xiommu1/oc8051_page_table_i/n956 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1469  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5] : \oc8051_xiommu1/oc8051_page_table_i/n957 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1470  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4] : \oc8051_xiommu1/oc8051_page_table_i/n958 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1471  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3] : \oc8051_xiommu1/oc8051_page_table_i/n959 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1472  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2] : \oc8051_xiommu1/oc8051_page_table_i/n960 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1473  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1] : \oc8051_xiommu1/oc8051_page_table_i/n961 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1474  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0] : \oc8051_xiommu1/oc8051_page_table_i/n962 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1475  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7] : \oc8051_xiommu1/oc8051_page_table_i/n963 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1476  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6] : \oc8051_xiommu1/oc8051_page_table_i/n964 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1477  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5] : \oc8051_xiommu1/oc8051_page_table_i/n965 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1478  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4] : \oc8051_xiommu1/oc8051_page_table_i/n966 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1479  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3] : \oc8051_xiommu1/oc8051_page_table_i/n967 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1480  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2] : \oc8051_xiommu1/oc8051_page_table_i/n968 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1481  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1] : \oc8051_xiommu1/oc8051_page_table_i/n969 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1482  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0] : \oc8051_xiommu1/oc8051_page_table_i/n970 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1483  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7] : \oc8051_xiommu1/oc8051_page_table_i/n971 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1484  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6] : \oc8051_xiommu1/oc8051_page_table_i/n972 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1485  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5] : \oc8051_xiommu1/oc8051_page_table_i/n973 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1486  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4] : \oc8051_xiommu1/oc8051_page_table_i/n974 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1487  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3] : \oc8051_xiommu1/oc8051_page_table_i/n975 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1488  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2] : \oc8051_xiommu1/oc8051_page_table_i/n976 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1489  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1] : \oc8051_xiommu1/oc8051_page_table_i/n977 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1490  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0] : \oc8051_xiommu1/oc8051_page_table_i/n978 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1491  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7] : \oc8051_xiommu1/oc8051_page_table_i/n979 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1492  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6] : \oc8051_xiommu1/oc8051_page_table_i/n980 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1493  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5] : \oc8051_xiommu1/oc8051_page_table_i/n981 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1494  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4] : \oc8051_xiommu1/oc8051_page_table_i/n982 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1495  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3] : \oc8051_xiommu1/oc8051_page_table_i/n983 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1496  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2] : \oc8051_xiommu1/oc8051_page_table_i/n984 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1497  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1] : \oc8051_xiommu1/oc8051_page_table_i/n985 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1498  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0] : \oc8051_xiommu1/oc8051_page_table_i/n986 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1499  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7] : \oc8051_xiommu1/oc8051_page_table_i/n987 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1500  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6] : \oc8051_xiommu1/oc8051_page_table_i/n988 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1501  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5] : \oc8051_xiommu1/oc8051_page_table_i/n989 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1502  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4] : \oc8051_xiommu1/oc8051_page_table_i/n990 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1503  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3] : \oc8051_xiommu1/oc8051_page_table_i/n991 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1504  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2] : \oc8051_xiommu1/oc8051_page_table_i/n992 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1505  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1] : \oc8051_xiommu1/oc8051_page_table_i/n993 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1506  = _cvpt_2211 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0] : \oc8051_xiommu1/oc8051_page_table_i/n994 ;   // oc8051_page_table.v(111)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1507  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n995 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1508  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n996 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1509  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n997 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1510  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n998 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1511  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n999 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1512  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1000 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1513  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1001 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1514  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1002 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1515  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1003 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1516  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1004 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1517  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1005 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1518  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1006 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1519  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1007 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1520  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1008 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1521  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1009 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1522  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1010 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1523  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1011 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1524  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1012 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1525  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1013 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1526  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1014 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1527  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1015 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1528  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1016 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1529  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1017 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1530  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1018 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1531  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1019 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1532  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1020 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1533  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1021 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1534  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1022 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1535  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1023 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1536  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1024 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1537  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1025 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1538  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1026 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1539  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1027 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1540  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1028 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1541  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1029 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1542  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1030 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1543  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1031 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1544  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1032 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1545  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1033 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1546  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1034 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1547  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1035 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1548  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1036 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1549  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1037 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1550  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1038 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1551  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1039 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1552  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1040 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1553  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1041 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1554  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1042 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1555  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1043 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1556  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1044 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1557  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1045 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1558  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1046 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1559  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1047 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1560  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1048 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1561  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1049 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1562  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1050 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1563  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1051 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1564  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1052 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1565  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1053 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1566  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1054 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1567  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1055 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1568  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1056 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1569  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1057 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1570  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1058 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1571  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1059 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1572  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1060 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1573  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1061 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1574  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1062 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1575  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1063 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1576  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1064 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1577  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1065 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1578  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1066 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1579  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1067 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1580  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1068 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1581  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1069 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1582  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1070 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1583  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1071 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1584  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1072 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1585  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1073 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1586  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1074 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1587  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1075 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1588  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1076 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1589  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1077 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1590  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1078 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1591  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1079 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1592  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1080 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1593  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1081 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1594  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1082 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1595  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1083 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1596  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1084 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1597  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1085 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1598  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1086 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1599  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1087 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1600  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1088 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1601  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1089 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1602  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1090 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1603  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1091 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1604  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1092 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1605  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1093 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1606  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1094 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1607  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1095 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1608  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1096 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1609  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1097 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1610  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1098 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1611  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1099 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1612  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1100 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1613  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1101 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1614  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1102 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1615  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1103 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1616  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1104 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1617  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1105 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1618  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1106 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1619  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1107 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1620  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1108 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1621  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1109 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1622  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1110 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1623  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1111 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1624  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1112 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1625  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1113 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1626  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1114 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1627  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1115 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1628  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1116 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1629  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1117 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1630  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1118 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1631  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1119 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1632  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1120 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1633  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1121 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1634  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1122 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1635  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1123 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1636  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1124 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1637  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1125 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1638  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1126 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1639  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1127 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1640  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1128 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1641  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1129 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1642  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1130 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1643  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1131 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1644  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1132 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1645  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1133 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1646  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1134 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1647  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1135 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1648  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1136 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1649  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1137 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1650  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1138 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1651  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1139 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1652  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1140 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1653  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1141 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1654  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1142 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1655  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1143 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1656  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1144 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1657  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1145 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1658  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1146 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1659  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1147 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1660  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1148 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1661  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1149 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1662  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1150 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1663  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1151 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1664  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1152 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1665  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1153 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1666  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1154 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1667  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1155 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1668  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1156 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1669  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1157 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1670  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1158 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1671  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1159 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1672  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1160 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1673  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1161 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1674  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1162 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1675  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1163 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1676  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1164 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1677  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1165 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1678  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1166 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1679  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1167 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1680  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1168 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1681  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1169 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1682  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1170 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1683  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1171 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1684  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1172 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1685  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1173 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1686  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1174 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1687  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1175 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1688  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1176 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1689  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1177 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1690  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1178 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1691  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1179 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1692  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1180 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1693  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1181 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1694  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1182 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1695  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1183 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1696  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1184 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1697  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1185 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1698  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1186 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1699  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1187 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1700  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1188 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1701  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1189 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1702  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1190 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1703  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1191 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1704  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1192 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1705  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1193 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1706  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1194 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1707  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1195 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1708  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1196 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1709  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1197 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1710  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1198 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1711  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1199 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1712  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1200 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1713  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1201 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1714  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1202 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1715  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1203 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1716  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1204 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1717  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1205 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1718  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1206 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1719  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1207 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1720  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1208 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1721  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1209 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1722  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1210 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1723  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1211 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1724  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1212 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1725  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1213 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1726  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1214 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1727  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1215 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1728  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1216 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1729  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1217 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1730  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1218 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1731  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1219 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1732  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1220 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1733  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1221 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1734  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1222 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1735  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1223 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1736  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1224 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1737  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1225 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1738  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1226 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1739  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1227 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1740  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1228 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1741  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1229 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1742  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1230 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1743  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1231 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1744  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1232 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1745  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1233 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1746  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1234 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1747  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1235 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1748  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1236 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1749  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1237 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1750  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1238 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1751  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1239 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1752  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1240 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1753  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1241 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1754  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1242 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1755  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1243 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1756  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1244 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1757  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1245 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1758  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1246 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1759  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1247 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1760  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1248 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1761  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1249 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1762  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1250 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1763  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1251 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1764  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1252 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1765  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1253 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1766  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1254 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1767  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1255 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1768  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1256 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1769  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1257 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1770  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1258 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1771  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1259 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1772  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1260 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1773  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1261 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1774  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1262 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1775  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1263 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1776  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1264 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1777  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1265 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1778  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1266 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1779  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1267 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1780  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1268 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1781  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1269 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1782  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1270 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1783  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1271 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1784  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1272 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1785  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1273 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1786  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1274 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1787  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1275 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1788  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1276 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1789  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1277 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1790  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1278 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1791  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1279 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1792  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1280 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1793  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1281 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1794  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1282 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1795  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1283 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1796  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1284 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1797  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1285 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1798  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1286 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1799  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1287 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1800  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1288 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1801  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1289 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1802  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1290 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1803  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1291 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1804  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1292 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1805  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1293 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1806  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1294 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1807  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1295 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1808  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1296 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1809  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1297 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1810  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1298 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1811  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1299 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1812  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1300 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1813  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1301 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1814  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1302 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1815  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1303 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1816  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1304 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1817  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1305 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1818  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1306 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1819  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1307 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1820  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1308 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1821  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1309 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1822  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1310 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1823  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1311 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1824  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1312 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1825  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1313 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1826  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1314 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1827  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1315 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1828  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1316 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1829  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1317 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1830  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1318 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1831  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1319 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1832  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1320 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1833  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1321 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1834  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1322 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1835  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1323 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1836  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1324 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1837  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1325 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1838  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1326 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1839  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1327 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1840  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1328 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1841  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1329 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1842  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1330 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1843  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1331 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1844  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1332 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1845  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1333 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1846  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1334 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1847  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1335 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1848  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1336 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1849  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1337 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1850  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1338 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1851  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1339 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1852  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1340 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1853  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1341 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1854  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1342 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1855  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1343 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1856  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1344 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1857  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1345 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1858  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1346 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1859  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1347 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1860  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1348 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1861  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1349 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1862  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1350 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1863  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1351 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1864  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1352 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1865  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1353 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1866  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1354 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1867  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1355 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1868  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1356 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1869  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1357 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1870  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1358 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1871  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1359 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1872  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1360 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1873  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1361 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1874  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1362 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1875  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1363 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1876  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1364 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1877  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1365 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1878  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1366 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1879  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1367 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1880  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1368 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1881  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1369 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1882  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1370 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1883  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1371 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1884  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1372 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1885  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1373 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1886  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1374 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1887  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1375 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1888  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1376 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1889  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1377 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1890  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1378 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1891  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1379 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1892  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1380 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1893  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1381 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1894  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1382 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1895  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1383 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1896  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1384 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1897  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1385 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1898  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1386 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1899  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1387 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1900  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1388 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1901  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1389 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1902  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1390 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1903  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1391 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1904  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1392 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1905  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1393 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1906  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1394 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1907  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1395 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1908  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1396 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1909  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1397 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1910  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1398 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1911  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1399 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1912  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1400 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1913  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1401 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1914  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1402 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1915  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1403 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1916  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1404 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1917  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1405 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1918  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1406 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1919  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1407 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1920  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1408 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1921  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1409 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1922  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1410 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1923  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1411 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1924  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1412 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1925  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1413 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1926  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1414 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1927  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1415 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1928  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1416 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1929  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1417 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1930  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1418 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1931  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1419 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1932  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1420 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1933  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1421 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1934  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1422 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1935  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1423 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1936  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1424 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1937  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1425 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1938  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1426 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1939  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1427 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1940  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1428 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1941  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1429 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1942  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1430 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1943  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1431 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1944  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1432 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1945  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1433 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1946  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1434 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1947  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1435 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1948  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1436 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1949  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1437 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1950  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1438 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1951  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1439 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1952  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1440 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1953  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1441 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1954  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1442 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1955  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1443 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1956  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1444 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1957  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1445 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1958  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1446 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1959  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1447 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1960  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1448 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1961  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1449 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1962  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1450 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1963  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1451 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1964  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1452 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1965  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1453 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1966  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1454 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1967  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1455 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1968  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1456 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1969  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1457 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1970  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1458 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1971  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1459 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1972  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1460 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1973  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1461 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1974  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1462 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1975  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1463 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1976  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1464 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1977  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1465 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1978  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1466 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1979  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1467 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1980  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1468 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1981  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1469 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1982  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1470 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1983  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1471 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1984  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1472 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1985  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1473 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1986  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1474 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1987  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1475 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1988  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1476 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1989  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1477 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1990  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1478 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1991  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1479 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1992  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1480 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1993  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1481 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1994  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1482 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1995  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1483 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1996  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1484 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1997  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1485 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1998  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1486 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n1999  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1487 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2000  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1488 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2001  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1489 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2002  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1490 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2003  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1491 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2004  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1492 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2005  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1493 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2006  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1494 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2007  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1495 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2008  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1496 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2009  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1497 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2010  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1498 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2011  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1499 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2012  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1500 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2013  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1501 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2014  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1502 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2015  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1503 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2016  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1504 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2017  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1505 ;   // oc8051_page_table.v(112)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2018  = _cvpt_914 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n1506 ;   // oc8051_page_table.v(112)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1958  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1508 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1959  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1509 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1960  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1510 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1961  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1511 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1962  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1512 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1963  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1513 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1964  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1514 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1965  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1515 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1966  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1516 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1967  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1517 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1968  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1518 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1969  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1519 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1970  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1520 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1971  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1521 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1972  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1522 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1973  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1523 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1974  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1524 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1975  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1525 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1976  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1526 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1977  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1527 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1978  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1528 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1979  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1529 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1980  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1530 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1981  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1531 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1982  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1532 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1983  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1533 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1984  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1534 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1985  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1535 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1986  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1536 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1987  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1537 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1988  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1538 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1989  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1539 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1990  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1540 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1991  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1541 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1992  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1542 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1993  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1543 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1994  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1544 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1995  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1545 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1996  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1546 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1997  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1547 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1998  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1548 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1999  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1549 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2000  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1550 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2001  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1551 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2002  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1552 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2003  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1553 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2004  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1554 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2005  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1555 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2006  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1556 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2007  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1557 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2008  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1558 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2009  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1559 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2010  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1560 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2011  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1561 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2012  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1562 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2013  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1563 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2014  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1564 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2015  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1565 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2016  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1566 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2017  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1567 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2018  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1568 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2019  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1569 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2020  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1570 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2021  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1571 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2022  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1572 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2023  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1573 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2024  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1574 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2025  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1575 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2026  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1576 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2027  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1577 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2028  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1578 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2029  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1579 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2030  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1580 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2031  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1581 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2032  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1582 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2033  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1583 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2034  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1584 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2035  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1585 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2036  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1586 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2037  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1587 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2038  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1588 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2039  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1589 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2040  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1590 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2041  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1591 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2042  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1592 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2043  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1593 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2044  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1594 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2045  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1595 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2046  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1596 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2047  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1597 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2048  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1598 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2049  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1599 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2050  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1600 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2051  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1601 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2052  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1602 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2053  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1603 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2054  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1604 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2055  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1605 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2056  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1606 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2057  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1607 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2058  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1608 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2059  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1609 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2060  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1610 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2061  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1611 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2062  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1612 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2063  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1613 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2064  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1614 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2065  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1615 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2066  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1616 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2067  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1617 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2068  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1618 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2069  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1619 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2070  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1620 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2071  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1621 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2072  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1622 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2073  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1623 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2074  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1624 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2075  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1625 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2076  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1626 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2077  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1627 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2078  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1628 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2079  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1629 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2080  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1630 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2081  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1631 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2082  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1632 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2083  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1633 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2084  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1634 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2085  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1635 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2086  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1636 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2087  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1637 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2088  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1638 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2089  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1639 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2090  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1640 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2091  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1641 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2092  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1642 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2093  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1643 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2094  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1644 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2095  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1645 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2096  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1646 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2097  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1647 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2098  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1648 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2099  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1649 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2100  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1650 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2101  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1651 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2102  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1652 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2103  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1653 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2104  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1654 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2105  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1655 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2106  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1656 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2107  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1657 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2108  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1658 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2109  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1659 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2110  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1660 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2111  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1661 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2112  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1662 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2113  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1663 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2114  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1664 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2115  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1665 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2116  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1666 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2117  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1667 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2118  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1668 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2119  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1669 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2120  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1670 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2121  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1671 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2122  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1672 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2123  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1673 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2124  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1674 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2125  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1675 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2126  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1676 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2127  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1677 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2128  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1678 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2129  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1679 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2130  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1680 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2131  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1681 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2132  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1682 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2133  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1683 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2134  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1684 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2135  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1685 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2136  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1686 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2137  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1687 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2138  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1688 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2139  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1689 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2140  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1690 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2141  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1691 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2142  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1692 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2143  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1693 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2144  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1694 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2145  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1695 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2146  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1696 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2147  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1697 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2148  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1698 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2149  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1699 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2150  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1700 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2151  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1701 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2152  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1702 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2153  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1703 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2154  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1704 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2155  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1705 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2156  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1706 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2157  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1707 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2158  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1708 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2159  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1709 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2160  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1710 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2161  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1711 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2162  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1712 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2163  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1713 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2164  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1714 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2165  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1715 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2166  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1716 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2167  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1717 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2168  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1718 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2169  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1719 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2170  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1720 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2171  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1721 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2172  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1722 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2173  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1723 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2174  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1724 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2175  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1725 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2176  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1726 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2177  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1727 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2178  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1728 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2179  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1729 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2180  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1730 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2181  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1731 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2182  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1732 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2183  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1733 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2184  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1734 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2185  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1735 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2186  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1736 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2187  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1737 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2188  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1738 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2189  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1739 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2190  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1740 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2191  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1741 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2192  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1742 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2193  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1743 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2194  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1744 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2195  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1745 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2196  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1746 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2197  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1747 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2198  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1748 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2199  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1749 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2200  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1750 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2201  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1751 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2202  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1752 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2203  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1753 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2204  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1754 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[1] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2205  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1755 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2206  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1756 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2207  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1757 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2208  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1758 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2209  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1759 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2210  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1760 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2211  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1761 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2212  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1762 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[0] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2213  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1763 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2214  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1764 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2215  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1765 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2216  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1766 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2217  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1767 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2218  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1768 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2219  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1769 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2220  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1770 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2221  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1771 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2222  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1772 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2223  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1773 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2224  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1774 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2225  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1775 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2226  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1776 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2227  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1777 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2228  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1778 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2229  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1779 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2230  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1780 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2231  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1781 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2232  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1782 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2233  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1783 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2234  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1784 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2235  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1785 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2236  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1786 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2237  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1787 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2238  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1788 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2239  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1789 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2240  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1790 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2241  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1791 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2242  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1792 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2243  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1793 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2244  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1794 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2245  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1795 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2246  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1796 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2247  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1797 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2248  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1798 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2249  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1799 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2250  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1800 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2251  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1801 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2252  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1802 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2253  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1803 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2254  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1804 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2255  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1805 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2256  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1806 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2257  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1807 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2258  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1808 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2259  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1809 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2260  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1810 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2261  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1811 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2262  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1812 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2263  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1813 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2264  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1814 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2265  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1815 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2266  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1816 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2267  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1817 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2268  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1818 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2269  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1819 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2270  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1820 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2271  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1821 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2272  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1822 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2273  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1823 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2274  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1824 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2275  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1825 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2276  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1826 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2277  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1827 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2278  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1828 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2279  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1829 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2280  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1830 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2281  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1831 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2282  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1832 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2283  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1833 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2284  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1834 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2285  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1835 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2286  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1836 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2287  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1837 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2288  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1838 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2289  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1839 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2290  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1840 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2291  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1841 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2292  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1842 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2293  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1843 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2294  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1844 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2295  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1845 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2296  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1846 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2297  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1847 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2298  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1848 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2299  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1849 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2300  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1850 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2301  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1851 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2302  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1852 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2303  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1853 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2304  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1854 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2305  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1855 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2306  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1856 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2307  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1857 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2308  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1858 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2309  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1859 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2310  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1860 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2311  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1861 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2312  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1862 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2313  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1863 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2314  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1864 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2315  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1865 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2316  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1866 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2317  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1867 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2318  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1868 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2319  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1869 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2320  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1870 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2321  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1871 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2322  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1872 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2323  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1873 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2324  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1874 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2325  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1875 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2326  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1876 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2327  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1877 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2328  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1878 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2329  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1879 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2330  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1880 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2331  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1881 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2332  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1882 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2333  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1883 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2334  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1884 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2335  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1885 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2336  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1886 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2337  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1887 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2338  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1888 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2339  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1889 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2340  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1890 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2341  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1891 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2342  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1892 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2343  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1893 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2344  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1894 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2345  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1895 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2346  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1896 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2347  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1897 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2348  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1898 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2349  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1899 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2350  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1900 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2351  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1901 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2352  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1902 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2353  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1903 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2354  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1904 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2355  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1905 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2356  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1906 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2357  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1907 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2358  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1908 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2359  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1909 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2360  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1910 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2361  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1911 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2362  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1912 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2363  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1913 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2364  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1914 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2365  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1915 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2366  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1916 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2367  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1917 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2368  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1918 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2369  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1919 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2370  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1920 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2371  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1921 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2372  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1922 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2373  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1923 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2374  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1924 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2375  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1925 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2376  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1926 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2377  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1927 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2378  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1928 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2379  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1929 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2380  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1930 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2381  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1931 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2382  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1932 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2383  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1933 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2384  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1934 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2385  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1935 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2386  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1936 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2387  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1937 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2388  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1938 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2389  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1939 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2390  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1940 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2391  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1941 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2392  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1942 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2393  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1943 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2394  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1944 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2395  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1945 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2396  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1946 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2397  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1947 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2398  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1948 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2399  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1949 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2400  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1950 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2401  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1951 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2402  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1952 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2403  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1953 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2404  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1954 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2405  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1955 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2406  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1956 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2407  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1957 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2408  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1958 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2409  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1959 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2410  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1960 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2411  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1961 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2412  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1962 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2413  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1963 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2414  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1964 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2415  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1965 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2416  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1966 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2417  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1967 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2418  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1968 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2419  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1969 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2420  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1970 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2421  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1971 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2422  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1972 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2423  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1973 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2424  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1974 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2425  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1975 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2426  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1976 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2427  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1977 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2428  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1978 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2429  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1979 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2430  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1980 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2431  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1981 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2432  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1982 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2433  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1983 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2434  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1984 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2435  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1985 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2436  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1986 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2437  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1987 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2438  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1988 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2439  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1989 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2440  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1990 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2441  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1991 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2442  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1992 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2443  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1993 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2444  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1994 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2445  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1995 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2446  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1996 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2447  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1997 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2448  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1998 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2449  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1999 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2450  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2000 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2451  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2001 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2452  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2002 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2453  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2003 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2454  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2004 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2455  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2005 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2456  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2006 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2457  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2007 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2458  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2008 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2459  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2009 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2460  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2010 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[1] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2461  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2011 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [7]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2462  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2012 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [6]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2463  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2013 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [5]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2464  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2014 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [4]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2465  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2015 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [3]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2466  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2016 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [2]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2467  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2017 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [1]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2468  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2018 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/rd_enabled[0] [0]));   // oc8051_page_table.v(113)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2607  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2632 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [15]));   // oc8051_page_table.v(169)
    and (\oc8051_xiommu1/oc8051_page_table_i/n2531 , \oc8051_xiommu1/stb_out , 
        \oc8051_xiommu1/wr_out ) ;   // oc8051_page_table.v(125)
    not (\oc8051_xiommu1/oc8051_page_table_i/n2532 , \oc8051_xiommu1/wr_en ) ;   // oc8051_page_table.v(125)
    and (_cvpt_3314, \oc8051_xiommu1/oc8051_page_table_i/n2531 , \oc8051_xiommu1/oc8051_page_table_i/n2532 ) ;   // oc8051_page_table.v(125)
    not (\oc8051_xiommu1/oc8051_page_table_i/n2534 , \oc8051_xiommu1/wr_out ) ;   // oc8051_page_table.v(126)
    and (\oc8051_xiommu1/oc8051_page_table_i/n2535 , \oc8051_xiommu1/stb_out , 
        \oc8051_xiommu1/oc8051_page_table_i/n2534 ) ;   // oc8051_page_table.v(126)
    not (\oc8051_xiommu1/oc8051_page_table_i/n2536 , \oc8051_xiommu1/rd_en ) ;   // oc8051_page_table.v(126)
    and (_cvpt_3312, \oc8051_xiommu1/oc8051_page_table_i/n2535 , \oc8051_xiommu1/oc8051_page_table_i/n2536 ) ;   // oc8051_page_table.v(126)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2542  = _cvpt_1209 ? \oc8051_xiommu1/selected_port [0] : 1'b1;   // oc8051_page_table.v(130)
    assign \oc8051_xiommu1/oc8051_page_table_i/accesser  = _cvpt_3236 ? \oc8051_xiommu1/selected_port [0] : \oc8051_xiommu1/oc8051_page_table_i/n2542 ;   // oc8051_page_table.v(130)
    or (_cvpt_3237, _cvpt_3314, _cvpt_3312) ;   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [15] = _cvpt_3237 ? _cvpt_3494 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [15];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [14] = _cvpt_3237 ? _cvpt_3478 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [14];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [13] = _cvpt_3237 ? _cvpt_3470 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [13];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [12] = _cvpt_3237 ? _cvpt_3466 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [12];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [11] = _cvpt_3237 ? _cvpt_1377 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [11];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [10] = _cvpt_3237 ? _cvpt_3710 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [10];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [9] = _cvpt_3237 ? _cvpt_3706 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [9];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [8] = _cvpt_3237 ? _cvpt_1401 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [8];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [7] = _cvpt_3237 ? \oc8051_xiommu1/addr_out [7] : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [7];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [6] = _cvpt_3237 ? \oc8051_xiommu1/addr_out [6] : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [6];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [5] = _cvpt_3237 ? \oc8051_xiommu1/addr_out [5] : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [5];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [4] = _cvpt_3237 ? _cvpt_3986 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [4];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [3] = _cvpt_3237 ? _cvpt_3970 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [3];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [2] = _cvpt_3237 ? _cvpt_3962 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [2];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [1] = _cvpt_3237 ? _cvpt_3958 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [1];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [0] = _cvpt_3237 ? _cvpt_1411 : \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [0];   // oc8051_page_table.v(132)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [2] = _cvpt_3237 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/illegal_src [2];   // oc8051_page_table.v(133)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [1] = _cvpt_3237 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/illegal_src [1];   // oc8051_page_table.v(133)
    assign \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [0] = _cvpt_3237 ? \oc8051_xiommu1/oc8051_page_table_i/accesser  : \oc8051_xiommu1/oc8051_page_table_i/illegal_src [0];   // oc8051_page_table.v(133)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2567  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [7] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [15];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2568  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [6] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [14];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2569  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [5] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [13];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2570  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [4] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [12];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2571  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [3] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [11];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2572  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [2] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [10];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2573  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [1] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [9];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2574  = _cvpt_3256 ? \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [0] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [8];   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2575  = _cvpt_3264 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2567 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2576  = _cvpt_3264 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2568 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2577  = _cvpt_3264 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2569 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2578  = _cvpt_3264 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2570 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2579  = _cvpt_3264 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2571 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2580  = _cvpt_3264 ? \oc8051_xiommu1/oc8051_page_table_i/illegal_src [2] : \oc8051_xiommu1/oc8051_page_table_i/n2572 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2581  = _cvpt_3264 ? \oc8051_xiommu1/oc8051_page_table_i/illegal_src [1] : \oc8051_xiommu1/oc8051_page_table_i/n2573 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2582  = _cvpt_3264 ? \oc8051_xiommu1/oc8051_page_table_i/illegal_src [0] : \oc8051_xiommu1/oc8051_page_table_i/n2574 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2583  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [15] : \oc8051_xiommu1/oc8051_page_table_i/n2575 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2584  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [14] : \oc8051_xiommu1/oc8051_page_table_i/n2576 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2585  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [13] : \oc8051_xiommu1/oc8051_page_table_i/n2577 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2586  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [12] : \oc8051_xiommu1/oc8051_page_table_i/n2578 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2587  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [11] : \oc8051_xiommu1/oc8051_page_table_i/n2579 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2588  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [10] : \oc8051_xiommu1/oc8051_page_table_i/n2580 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2589  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [9] : \oc8051_xiommu1/oc8051_page_table_i/n2581 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2590  = _cvpt_3272 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [8] : \oc8051_xiommu1/oc8051_page_table_i/n2582 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2591  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [7] : \oc8051_xiommu1/oc8051_page_table_i/n2583 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2592  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [6] : \oc8051_xiommu1/oc8051_page_table_i/n2584 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2593  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [5] : \oc8051_xiommu1/oc8051_page_table_i/n2585 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2594  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [4] : \oc8051_xiommu1/oc8051_page_table_i/n2586 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2595  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [3] : \oc8051_xiommu1/oc8051_page_table_i/n2587 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2596  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [2] : \oc8051_xiommu1/oc8051_page_table_i/n2588 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2597  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [1] : \oc8051_xiommu1/oc8051_page_table_i/n2589 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2598  = _cvpt_3280 ? \oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [0] : \oc8051_xiommu1/oc8051_page_table_i/n2590 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [7] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2591 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [6] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2592 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [5] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2593 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [4] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2594 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [3] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2595 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [2] = _cvpt_3288 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2596 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [1] = _cvpt_3288 ? \oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [1] : \oc8051_xiommu1/oc8051_page_table_i/n2597 ;   // oc8051_page_table.v(139)
    assign \oc8051_xiommu1/data_out_ia [0] = _cvpt_3288 ? \oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [0] : \oc8051_xiommu1/oc8051_page_table_i/n2598 ;   // oc8051_page_table.v(139)
    and (\oc8051_xiommu1/ack_ia , _cvpt_111, \oc8051_xiommu1/ia_addr_range ) ;   // oc8051_page_table.v(141)
    not (\oc8051_xiommu1/oc8051_page_table_i/n2610 , \oc8051_xiommu1/oc8051_page_table_i/accesser ) ;   // oc8051_page_table.v(157)
    and (_cvpt_3296, _cvpt_3237, \oc8051_xiommu1/oc8051_page_table_i/n2610 ) ;   // oc8051_page_table.v(157)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2612  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [15] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [15];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2613  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [14] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [14];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2614  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [13] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [13];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2615  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [12] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [12];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2616  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [11] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [11];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2617  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [10] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [10];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2618  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [9] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [9];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2619  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [8] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [8];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2620  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [7] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [7];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2621  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [6] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [6];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2622  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [5] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [5];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2623  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [4] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [4];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2624  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [3] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [3];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2625  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [2] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [2];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2626  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [1] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [1];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2627  = _cvpt_3296 ? \oc8051_xiommu1/dpc_ot [0] : \oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [0];   // oc8051_page_table.v(159)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2628  = _cvpt_3312 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [1];   // oc8051_page_table.v(167)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2629  = _cvpt_3312 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [0];   // oc8051_page_table.v(167)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2630  = _cvpt_3314 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2628 ;   // oc8051_page_table.v(167)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2631  = _cvpt_3314 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/n2629 ;   // oc8051_page_table.v(167)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2632  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [15];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2633  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [14];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2634  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [13];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2635  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [12];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2636  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [11];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2637  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [10];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2638  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [9];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2639  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [8];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2640  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [7];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2641  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [6];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2642  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [5];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2643  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [4];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2644  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [3];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2645  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [2];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2646  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [1];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2647  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_reg_next [0];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2648  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2630 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2649  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2631 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2650  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [2];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2651  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [1];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2652  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/ia_src_next [0];   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2653  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2612 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2654  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2613 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2655  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2614 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2656  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2615 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2657  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2616 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2658  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2617 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2659  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2618 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2660  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2619 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2661  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2620 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2662  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2621 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2663  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2622 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2664  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2623 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2665  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2624 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2666  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2625 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2667  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2626 ;   // oc8051_page_table.v(168)
    assign \oc8051_xiommu1/oc8051_page_table_i/n2668  = _cvpt_914 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/n2627 ;   // oc8051_page_table.v(168)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2608  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2633 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [14]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2609  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2634 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [13]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2610  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2635 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [12]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2611  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2636 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [11]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2612  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2637 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [10]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2613  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2638 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [9]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2614  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2639 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [8]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2615  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2640 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [7]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2616  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2641 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [6]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2617  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2642 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [5]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2618  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2643 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [4]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2619  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2644 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [3]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2620  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2645 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [2]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2621  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2646 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [1]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2622  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2647 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_addr_reg [0]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2623  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2648 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [1]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2624  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2649 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/ia_rwn_reg [0]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2625  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2650 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/illegal_src [2]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2626  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2651 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/illegal_src [1]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2627  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2652 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/illegal_src [0]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2628  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2653 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [15]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2629  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2654 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [14]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2630  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2655 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [13]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2631  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2656 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [12]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2632  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2657 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [11]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2633  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2658 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [10]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2634  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2659 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [9]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2635  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2660 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [8]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2636  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2661 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [7]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2637  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2662 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [6]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2638  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2663 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [5]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2639  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2664 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [4]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2640  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2665 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [3]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2641  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2666 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [2]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2642  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2667 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [1]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i2643  (.d(\oc8051_xiommu1/oc8051_page_table_i/n2668 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/pc_ia_reg [0]));   // oc8051_page_table.v(169)
    VERIFIC_DFFRS \oc8051_xiommu1/oc8051_page_table_i/i1957  (.d(\oc8051_xiommu1/oc8051_page_table_i/n1507 ), 
            .clk(clk), .s(1'b0), .r(1'b0), .q(\oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [7]));   // oc8051_page_table.v(113)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n2  = _cvpt_3353 ? \oc8051_xiommu1/proc_addr [0] : 1'b1;   // aes_top.v(94)
    xor (_cvpt_3354, 1'b0, \oc8051_xiommu1/proc_addr [1]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n4  = _cvpt_3354 ? \oc8051_xiommu1/proc_addr [1] : \oc8051_xiommu1/aes_top_i/LessThan_3/n2 ;   // aes_top.v(94)
    xor (_cvpt_3355, 1'b0, \oc8051_xiommu1/proc_addr [2]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n6  = _cvpt_3355 ? \oc8051_xiommu1/proc_addr [2] : \oc8051_xiommu1/aes_top_i/LessThan_3/n4 ;   // aes_top.v(94)
    xor (_cvpt_3356, 1'b0, \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n8  = _cvpt_3356 ? \oc8051_xiommu1/proc_addr [3] : \oc8051_xiommu1/aes_top_i/LessThan_3/n6 ;   // aes_top.v(94)
    xor (_cvpt_3357, 1'b0, \oc8051_xiommu1/proc_addr [4]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n10  = _cvpt_3357 ? \oc8051_xiommu1/proc_addr [4] : \oc8051_xiommu1/aes_top_i/LessThan_3/n8 ;   // aes_top.v(94)
    xor (_cvpt_3358, 1'b0, \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n12  = _cvpt_3358 ? \oc8051_xiommu1/proc_addr [5] : \oc8051_xiommu1/aes_top_i/LessThan_3/n10 ;   // aes_top.v(94)
    xor (_cvpt_3359, 1'b0, \oc8051_xiommu1/proc_addr [6]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n14  = _cvpt_3359 ? \oc8051_xiommu1/proc_addr [6] : \oc8051_xiommu1/aes_top_i/LessThan_3/n12 ;   // aes_top.v(94)
    xor (_cvpt_3360, 1'b0, \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n16  = _cvpt_3360 ? \oc8051_xiommu1/proc_addr [7] : \oc8051_xiommu1/aes_top_i/LessThan_3/n14 ;   // aes_top.v(94)
    xor (_cvpt_3361, 1'b1, \oc8051_xiommu1/proc_addr [8]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n18  = _cvpt_3361 ? \oc8051_xiommu1/proc_addr [8] : \oc8051_xiommu1/aes_top_i/LessThan_3/n16 ;   // aes_top.v(94)
    xor (_cvpt_3362, 1'b1, \oc8051_xiommu1/proc_addr [9]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n20  = _cvpt_3362 ? \oc8051_xiommu1/proc_addr [9] : \oc8051_xiommu1/aes_top_i/LessThan_3/n18 ;   // aes_top.v(94)
    xor (_cvpt_3363, 1'b1, \oc8051_xiommu1/proc_addr [10]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n22  = _cvpt_3363 ? \oc8051_xiommu1/proc_addr [10] : \oc8051_xiommu1/aes_top_i/LessThan_3/n20 ;   // aes_top.v(94)
    xor (_cvpt_3364, 1'b1, \oc8051_xiommu1/proc_addr [11]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n24  = _cvpt_3364 ? \oc8051_xiommu1/proc_addr [11] : \oc8051_xiommu1/aes_top_i/LessThan_3/n22 ;   // aes_top.v(94)
    xor (_cvpt_3365, 1'b1, \oc8051_xiommu1/proc_addr [12]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n26  = _cvpt_3365 ? \oc8051_xiommu1/proc_addr [12] : \oc8051_xiommu1/aes_top_i/LessThan_3/n24 ;   // aes_top.v(94)
    xor (_cvpt_3366, 1'b1, \oc8051_xiommu1/proc_addr [13]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n28  = _cvpt_3366 ? \oc8051_xiommu1/proc_addr [13] : \oc8051_xiommu1/aes_top_i/LessThan_3/n26 ;   // aes_top.v(94)
    xor (_cvpt_3367, 1'b1, \oc8051_xiommu1/proc_addr [14]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_3/n30  = _cvpt_3367 ? \oc8051_xiommu1/proc_addr [14] : \oc8051_xiommu1/aes_top_i/LessThan_3/n28 ;   // aes_top.v(94)
    xor (_cvpt_3368, 1'b1, \oc8051_xiommu1/proc_addr [15]) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/n4  = _cvpt_3368 ? \oc8051_xiommu1/proc_addr [15] : \oc8051_xiommu1/aes_top_i/LessThan_3/n30 ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n2  = _cvpt_3369 ? 1'b0 : 1'b0;   // aes_top.v(94)
    xor (_cvpt_3370, \oc8051_xiommu1/proc_addr [1], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n4  = _cvpt_3370 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n2 ;   // aes_top.v(94)
    xor (_cvpt_3371, \oc8051_xiommu1/proc_addr [2], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n6  = _cvpt_3371 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n4 ;   // aes_top.v(94)
    xor (_cvpt_3372, \oc8051_xiommu1/proc_addr [3], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n8  = _cvpt_3372 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n6 ;   // aes_top.v(94)
    xor (_cvpt_3373, \oc8051_xiommu1/proc_addr [4], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n10  = _cvpt_3373 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n8 ;   // aes_top.v(94)
    xor (_cvpt_3374, \oc8051_xiommu1/proc_addr [5], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n12  = _cvpt_3374 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n10 ;   // aes_top.v(94)
    xor (_cvpt_3375, \oc8051_xiommu1/proc_addr [6], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n14  = _cvpt_3375 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n12 ;   // aes_top.v(94)
    xor (_cvpt_3376, \oc8051_xiommu1/proc_addr [7], 1'b0) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n16  = _cvpt_3376 ? 1'b0 : \oc8051_xiommu1/aes_top_i/LessThan_4/n14 ;   // aes_top.v(94)
    xor (_cvpt_3377, \oc8051_xiommu1/proc_addr [8], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n18  = _cvpt_3377 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n16 ;   // aes_top.v(94)
    xor (_cvpt_3378, \oc8051_xiommu1/proc_addr [9], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n20  = _cvpt_3378 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n18 ;   // aes_top.v(94)
    xor (_cvpt_3379, \oc8051_xiommu1/proc_addr [10], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n22  = _cvpt_3379 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n20 ;   // aes_top.v(94)
    xor (_cvpt_3380, \oc8051_xiommu1/proc_addr [11], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n24  = _cvpt_3380 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n22 ;   // aes_top.v(94)
    xor (_cvpt_3381, \oc8051_xiommu1/proc_addr [12], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n26  = _cvpt_3381 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n24 ;   // aes_top.v(94)
    xor (_cvpt_3382, \oc8051_xiommu1/proc_addr [13], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n28  = _cvpt_3382 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n26 ;   // aes_top.v(94)
    xor (_cvpt_3383, \oc8051_xiommu1/proc_addr [14], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/LessThan_4/n30  = _cvpt_3383 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n28 ;   // aes_top.v(94)
    xor (_cvpt_3384, \oc8051_xiommu1/proc_addr [15], 1'b1) ;   // aes_top.v(94)
    assign \oc8051_xiommu1/aes_top_i/n5  = _cvpt_3384 ? 1'b1 : \oc8051_xiommu1/aes_top_i/LessThan_4/n30 ;   // aes_top.v(94)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n2 , \oc8051_xiommu1/proc_addr [2], 
        \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n2 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n4 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n5 , \oc8051_xiommu1/proc_addr [6], 
        \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n5 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n6 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n8 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n9 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/n11 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n9 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n11 , \oc8051_xiommu1/aes_top_i/n12 , 
        \oc8051_xiommu1/aes_top_i/n13 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n12 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n12 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n13 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_15/n15 , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_15/n14 ) ;   // aes_top.v(97)
    not (\oc8051_xiommu1/aes_top_i/sel_reg_start , \oc8051_xiommu1/aes_top_i/reduce_nor_15/n15 ) ;   // aes_top.v(97)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n2 , \oc8051_xiommu1/proc_addr [2], 
        \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n2 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n4 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n5 , \oc8051_xiommu1/proc_addr [6], 
        \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n5 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n6 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n8 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n9 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/n11 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n9 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n11 , \oc8051_xiommu1/aes_top_i/n12 , 
        \oc8051_xiommu1/aes_top_i/n13 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n12 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n12 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n13 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_25/n15 , \oc8051_xiommu1/aes_top_i/reduce_nor_25/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_25/n14 ) ;   // aes_top.v(98)
    not (_cvpt_327, \oc8051_xiommu1/aes_top_i/reduce_nor_25/n15 ) ;   // aes_top.v(98)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n2 , \oc8051_xiommu1/aes_top_i/n28 , 
        \oc8051_xiommu1/proc_addr [3]) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n2 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n4 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n5 , \oc8051_xiommu1/proc_addr [6], 
        \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n4 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n5 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n7 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n6 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n8 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n9 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/n11 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n8 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n9 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n11 , \oc8051_xiommu1/aes_top_i/n12 , 
        \oc8051_xiommu1/aes_top_i/n13 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n12 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n11 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n12 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n13 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_36/n15 , \oc8051_xiommu1/aes_top_i/reduce_nor_36/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_36/n14 ) ;   // aes_top.v(99)
    not (_cvpt_303, \oc8051_xiommu1/aes_top_i/reduce_nor_36/n15 ) ;   // aes_top.v(99)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n2 , \oc8051_xiommu1/aes_top_i/n27 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n1 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n3 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n4 , \oc8051_xiommu1/proc_addr [6], 
        \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n4 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n5 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n7 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n8 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/n11 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n8 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n10 , \oc8051_xiommu1/aes_top_i/n12 , 
        \oc8051_xiommu1/aes_top_i/n13 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n11 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n12 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n11 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n9 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n12 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_46/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_46/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_46/n13 ) ;   // aes_top.v(100)
    not (_cvpt_319, \oc8051_xiommu1/aes_top_i/reduce_nor_46/n14 ) ;   // aes_top.v(100)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n2 , \oc8051_xiommu1/proc_addr [1], 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n1 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n3 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/proc_addr [5]) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n4 , \oc8051_xiommu1/proc_addr [6], 
        \oc8051_xiommu1/proc_addr [7]) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n3 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n4 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n6 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n5 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n7 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n8 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/n11 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n9 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n8 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n10 , \oc8051_xiommu1/aes_top_i/n12 , 
        \oc8051_xiommu1/aes_top_i/n13 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n11 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n12 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n11 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n13 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n9 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n12 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_56/n14 , \oc8051_xiommu1/aes_top_i/reduce_nor_56/n6 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_56/n13 ) ;   // aes_top.v(101)
    not (_cvpt_311, \oc8051_xiommu1/aes_top_i/reduce_nor_56/n14 ) ;   // aes_top.v(101)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n2 , \oc8051_xiommu1/aes_top_i/n58 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n1 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n3 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n4 , \oc8051_xiommu1/proc_addr [7], 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n3 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n4 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n6 , \oc8051_xiommu1/aes_top_i/n11 , 
        \oc8051_xiommu1/aes_top_i/n12 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n7 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n6 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n8 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n9 , \oc8051_xiommu1/aes_top_i/n13 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n8 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n9 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_66/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_66/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_66/n10 ) ;   // aes_top.v(102)
    not (_cvpt_295, \oc8051_xiommu1/aes_top_i/reduce_nor_66/n11 ) ;   // aes_top.v(102)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n2 , \oc8051_xiommu1/proc_addr [4], 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n1 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n3 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n4 , \oc8051_xiommu1/proc_addr [7], 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n3 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n4 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n6 , \oc8051_xiommu1/aes_top_i/n11 , 
        \oc8051_xiommu1/aes_top_i/n12 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n7 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n6 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n8 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n9 , \oc8051_xiommu1/aes_top_i/n13 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n8 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n9 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_76/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_76/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_76/n10 ) ;   // aes_top.v(103)
    not (_cvpt_287, \oc8051_xiommu1/aes_top_i/reduce_nor_76/n11 ) ;   // aes_top.v(103)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n2 , \oc8051_xiommu1/aes_top_i/n58 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n1 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n3 , \oc8051_xiommu1/aes_top_i/n8 , 
        \oc8051_xiommu1/aes_top_i/n9 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n4 , \oc8051_xiommu1/proc_addr [7], 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n3 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n5 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n2 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n4 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n6 , \oc8051_xiommu1/aes_top_i/n11 , 
        \oc8051_xiommu1/aes_top_i/n12 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n7 , \oc8051_xiommu1/aes_top_i/n10 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n6 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n8 , \oc8051_xiommu1/aes_top_i/n14 , 
        \oc8051_xiommu1/aes_top_i/n15 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n9 , \oc8051_xiommu1/aes_top_i/n13 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n8 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n10 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n7 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n9 ) ;   // aes_top.v(104)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_87/n11 , \oc8051_xiommu1/aes_top_i/reduce_nor_87/n5 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_87/n10 ) ;   // aes_top.v(104)
    not (_cvpt_279, \oc8051_xiommu1/aes_top_i/reduce_nor_87/n11 ) ;   // aes_top.v(104)
    not (_cvpt_408, \oc8051_xiommu1/aes_top_i/reduce_nor_144/n1 ) ;   // aes_top.v(120)
    not (_cvpt_406, \oc8051_xiommu1/aes_top_i/reduce_nor_146/n1 ) ;   // aes_top.v(121)
    not (_cvpt_404, \oc8051_xiommu1/aes_top_i/reduce_nor_148/n1 ) ;   // aes_top.v(122)
    not (_cvpt_402, \oc8051_xiommu1/aes_top_i/reduce_nor_151/n1 ) ;   // aes_top.v(123)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n2 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [5]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n175 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n4 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n4 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [6]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n174 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n6 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n6 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [7]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n173 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n8 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i5  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n8 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [8]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n172 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n10 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i6  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n10 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [9]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n171 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n12 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i7  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n12 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [10]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n170 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n14 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i8  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n14 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [11]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n169 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n16 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i9  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n16 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [12]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n168 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n18 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i10  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n18 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [13]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n167 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n20 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i11  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n20 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [14]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n166 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/n22 ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_163/i12  (.cin(\oc8051_xiommu1/aes_top_i/add_163/n22 ), 
            .a(\oc8051_xiommu1/aes_top_i/operated_bytes_count [15]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n165 ), .cout(\oc8051_xiommu1/aes_top_i/add_163/cout ));   // aes_top.v(214)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n2 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [5]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n218 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_194/n4 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n4 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [6]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n217 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_194/n6 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n6 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [7]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n216 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_194/n8 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i5  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n8 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [8]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n215 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_194/n10 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i6  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n10 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [9]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n214 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_194/n12 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i7  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n12 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [10]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n213 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n14 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i8  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n14 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [11]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n212 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n16 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i9  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n16 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [12]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n211 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n18 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i10  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n18 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [13]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n210 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n20 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i11  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n20 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [14]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n209 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/n22 ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_194/i12  (.cin(\oc8051_xiommu1/aes_top_i/add_194/n22 ), 
            .a(\oc8051_xiommu1/aes_top_i/block_counter [15]), .b(1'b0), 
            .o(\oc8051_xiommu1/aes_top_i/n208 ), .cout(\oc8051_xiommu1/aes_top_i/add_194/cout ));   // aes_top.v(220)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_225/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_225/n2 ), 
            .a(\oc8051_xiommu1/aes_top_i/byte_counter [1]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n253 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_225/n4 ));   // aes_top.v(228)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_225/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_225/n4 ), 
            .a(\oc8051_xiommu1/aes_top_i/byte_counter [2]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n252 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_225/n6 ));   // aes_top.v(228)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_225/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_225/n6 ), 
            .a(\oc8051_xiommu1/aes_top_i/byte_counter [3]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/n251 ), 
            .cout(\oc8051_xiommu1/aes_top_i/add_225/cout ));   // aes_top.v(228)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_240/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(231)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_240/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_240/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_240/n2 ) ;   // aes_top.v(231)
    not (\oc8051_xiommu1/aes_top_i/n269 , \oc8051_xiommu1/aes_top_i/reduce_nor_240/n3 ) ;   // aes_top.v(231)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n2  = _cvpt_3385 ? \oc8051_xiommu1/aes_len [0] : 1'b0;   // aes_top.v(234)
    xor (_cvpt_3386, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [1], 
        \oc8051_xiommu1/aes_len [1]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n4  = _cvpt_3386 ? \oc8051_xiommu1/aes_len [1] : \oc8051_xiommu1/aes_top_i/LessThan_243/n2 ;   // aes_top.v(234)
    xor (_cvpt_3387, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [2], 
        \oc8051_xiommu1/aes_len [2]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n6  = _cvpt_3387 ? \oc8051_xiommu1/aes_len [2] : \oc8051_xiommu1/aes_top_i/LessThan_243/n4 ;   // aes_top.v(234)
    xor (_cvpt_3388, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [3], 
        \oc8051_xiommu1/aes_len [3]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n8  = _cvpt_3388 ? \oc8051_xiommu1/aes_len [3] : \oc8051_xiommu1/aes_top_i/LessThan_243/n6 ;   // aes_top.v(234)
    xor (_cvpt_3389, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [4], 
        \oc8051_xiommu1/aes_len [4]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n10  = _cvpt_3389 ? \oc8051_xiommu1/aes_len [4] : \oc8051_xiommu1/aes_top_i/LessThan_243/n8 ;   // aes_top.v(234)
    xor (_cvpt_3390, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [5], 
        \oc8051_xiommu1/aes_len [5]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n12  = _cvpt_3390 ? \oc8051_xiommu1/aes_len [5] : \oc8051_xiommu1/aes_top_i/LessThan_243/n10 ;   // aes_top.v(234)
    xor (_cvpt_3391, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [6], 
        \oc8051_xiommu1/aes_len [6]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n14  = _cvpt_3391 ? \oc8051_xiommu1/aes_len [6] : \oc8051_xiommu1/aes_top_i/LessThan_243/n12 ;   // aes_top.v(234)
    xor (_cvpt_3392, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [7], 
        \oc8051_xiommu1/aes_len [7]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n16  = _cvpt_3392 ? \oc8051_xiommu1/aes_len [7] : \oc8051_xiommu1/aes_top_i/LessThan_243/n14 ;   // aes_top.v(234)
    xor (_cvpt_3393, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [8], 
        \oc8051_xiommu1/aes_len [8]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n18  = _cvpt_3393 ? \oc8051_xiommu1/aes_len [8] : \oc8051_xiommu1/aes_top_i/LessThan_243/n16 ;   // aes_top.v(234)
    xor (_cvpt_3394, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [9], 
        \oc8051_xiommu1/aes_len [9]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n20  = _cvpt_3394 ? \oc8051_xiommu1/aes_len [9] : \oc8051_xiommu1/aes_top_i/LessThan_243/n18 ;   // aes_top.v(234)
    xor (_cvpt_3395, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [10], 
        \oc8051_xiommu1/aes_len [10]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n22  = _cvpt_3395 ? \oc8051_xiommu1/aes_len [10] : \oc8051_xiommu1/aes_top_i/LessThan_243/n20 ;   // aes_top.v(234)
    xor (_cvpt_3396, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [11], 
        \oc8051_xiommu1/aes_len [11]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n24  = _cvpt_3396 ? \oc8051_xiommu1/aes_len [11] : \oc8051_xiommu1/aes_top_i/LessThan_243/n22 ;   // aes_top.v(234)
    xor (_cvpt_3397, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [12], 
        \oc8051_xiommu1/aes_len [12]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n26  = _cvpt_3397 ? \oc8051_xiommu1/aes_len [12] : \oc8051_xiommu1/aes_top_i/LessThan_243/n24 ;   // aes_top.v(234)
    xor (_cvpt_3398, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [13], 
        \oc8051_xiommu1/aes_len [13]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n28  = _cvpt_3398 ? \oc8051_xiommu1/aes_len [13] : \oc8051_xiommu1/aes_top_i/LessThan_243/n26 ;   // aes_top.v(234)
    xor (_cvpt_3399, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [14], 
        \oc8051_xiommu1/aes_len [14]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/LessThan_243/n30  = _cvpt_3399 ? \oc8051_xiommu1/aes_len [14] : \oc8051_xiommu1/aes_top_i/LessThan_243/n28 ;   // aes_top.v(234)
    xor (_cvpt_3400, \oc8051_xiommu1/aes_top_i/operated_bytes_count_next [15], 
        \oc8051_xiommu1/aes_len [15]) ;   // aes_top.v(234)
    assign \oc8051_xiommu1/aes_top_i/n272  = _cvpt_3400 ? \oc8051_xiommu1/aes_len [15] : \oc8051_xiommu1/aes_top_i/LessThan_243/n30 ;   // aes_top.v(234)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n2 ), 
            .a(\oc8051_xiommu1/aes_addr [1]), .b(\oc8051_xiommu1/aes_top_i/block_counter [1]), 
            .o(\oc8051_xiommu1/aes_top_i/n289 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n4 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n4 ), 
            .a(\oc8051_xiommu1/aes_addr [2]), .b(\oc8051_xiommu1/aes_top_i/block_counter [2]), 
            .o(\oc8051_xiommu1/aes_top_i/n288 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n6 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n6 ), 
            .a(\oc8051_xiommu1/aes_addr [3]), .b(\oc8051_xiommu1/aes_top_i/block_counter [3]), 
            .o(\oc8051_xiommu1/aes_top_i/n287 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n8 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i5  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n8 ), 
            .a(\oc8051_xiommu1/aes_addr [4]), .b(\oc8051_xiommu1/aes_top_i/block_counter [4]), 
            .o(\oc8051_xiommu1/aes_top_i/n286 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n10 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i6  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n10 ), 
            .a(\oc8051_xiommu1/aes_addr [5]), .b(\oc8051_xiommu1/aes_top_i/block_counter [5]), 
            .o(\oc8051_xiommu1/aes_top_i/n285 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n12 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i7  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n12 ), 
            .a(\oc8051_xiommu1/aes_addr [6]), .b(\oc8051_xiommu1/aes_top_i/block_counter [6]), 
            .o(\oc8051_xiommu1/aes_top_i/n284 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n14 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i8  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n14 ), 
            .a(\oc8051_xiommu1/aes_addr [7]), .b(\oc8051_xiommu1/aes_top_i/block_counter [7]), 
            .o(\oc8051_xiommu1/aes_top_i/n283 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n16 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i9  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n16 ), 
            .a(\oc8051_xiommu1/aes_addr [8]), .b(\oc8051_xiommu1/aes_top_i/block_counter [8]), 
            .o(\oc8051_xiommu1/aes_top_i/n282 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n18 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i10  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n18 ), 
            .a(\oc8051_xiommu1/aes_addr [9]), .b(\oc8051_xiommu1/aes_top_i/block_counter [9]), 
            .o(\oc8051_xiommu1/aes_top_i/n281 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n20 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i11  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n20 ), 
            .a(\oc8051_xiommu1/aes_addr [10]), .b(\oc8051_xiommu1/aes_top_i/block_counter [10]), 
            .o(\oc8051_xiommu1/aes_top_i/n280 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n22 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i12  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n22 ), 
            .a(\oc8051_xiommu1/aes_addr [11]), .b(\oc8051_xiommu1/aes_top_i/block_counter [11]), 
            .o(\oc8051_xiommu1/aes_top_i/n279 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n24 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i13  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n24 ), 
            .a(\oc8051_xiommu1/aes_addr [12]), .b(\oc8051_xiommu1/aes_top_i/block_counter [12]), 
            .o(\oc8051_xiommu1/aes_top_i/n278 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n26 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i14  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n26 ), 
            .a(\oc8051_xiommu1/aes_addr [13]), .b(\oc8051_xiommu1/aes_top_i/block_counter [13]), 
            .o(\oc8051_xiommu1/aes_top_i/n277 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n28 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i15  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n28 ), 
            .a(\oc8051_xiommu1/aes_addr [14]), .b(\oc8051_xiommu1/aes_top_i/block_counter [14]), 
            .o(\oc8051_xiommu1/aes_top_i/n276 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/n30 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_245/i16  (.cin(\oc8051_xiommu1/aes_top_i/add_245/n30 ), 
            .a(\oc8051_xiommu1/aes_addr [15]), .b(\oc8051_xiommu1/aes_top_i/block_counter [15]), 
            .o(\oc8051_xiommu1/aes_top_i/n275 ), .cout(\oc8051_xiommu1/aes_top_i/add_245/cout ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n2 ), 
            .a(\oc8051_xiommu1/aes_top_i/n289 ), .b(\oc8051_xiommu1/aes_top_i/byte_counter [1]), 
            .o(\oc8051_xiommu1/aes_xram_addr [1]), .cout(\oc8051_xiommu1/aes_top_i/add_246/n4 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n4 ), 
            .a(\oc8051_xiommu1/aes_top_i/n288 ), .b(\oc8051_xiommu1/aes_top_i/byte_counter [2]), 
            .o(\oc8051_xiommu1/aes_xram_addr [2]), .cout(\oc8051_xiommu1/aes_top_i/add_246/n6 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n6 ), 
            .a(\oc8051_xiommu1/aes_top_i/n287 ), .b(\oc8051_xiommu1/aes_top_i/byte_counter [3]), 
            .o(\oc8051_xiommu1/aes_xram_addr [3]), .cout(\oc8051_xiommu1/aes_top_i/add_246/n8 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i5  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n8 ), 
            .a(\oc8051_xiommu1/aes_top_i/n286 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [4]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n10 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i6  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n10 ), 
            .a(\oc8051_xiommu1/aes_top_i/n285 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [5]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n12 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i7  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n12 ), 
            .a(\oc8051_xiommu1/aes_top_i/n284 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [6]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n14 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i8  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n14 ), 
            .a(\oc8051_xiommu1/aes_top_i/n283 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [7]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n16 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i9  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n16 ), 
            .a(\oc8051_xiommu1/aes_top_i/n282 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [8]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n18 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i10  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n18 ), 
            .a(\oc8051_xiommu1/aes_top_i/n281 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [9]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n20 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i11  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n20 ), 
            .a(\oc8051_xiommu1/aes_top_i/n280 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [10]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n22 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i12  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n22 ), 
            .a(\oc8051_xiommu1/aes_top_i/n279 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [11]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n24 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i13  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n24 ), 
            .a(\oc8051_xiommu1/aes_top_i/n278 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [12]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n26 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i14  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n26 ), 
            .a(\oc8051_xiommu1/aes_top_i/n277 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [13]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n28 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i15  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n28 ), 
            .a(\oc8051_xiommu1/aes_top_i/n276 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [14]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/n30 ));   // aes_top.v(237)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_246/i16  (.cin(\oc8051_xiommu1/aes_top_i/add_246/n30 ), 
            .a(\oc8051_xiommu1/aes_top_i/n275 ), .b(1'b0), .o(\oc8051_xiommu1/aes_xram_addr [15]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_246/cout ));   // aes_top.v(237)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_265/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(263)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_265/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_265/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_265/n2 ) ;   // aes_top.v(263)
    not (_cvpt_906, \oc8051_xiommu1/aes_top_i/reduce_nor_265/n3 ) ;   // aes_top.v(263)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_276/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(264)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_276/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_276/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_276/n2 ) ;   // aes_top.v(264)
    not (_cvpt_898, \oc8051_xiommu1/aes_top_i/reduce_nor_276/n3 ) ;   // aes_top.v(264)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_287/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(265)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_287/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_287/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_287/n2 ) ;   // aes_top.v(265)
    not (_cvpt_890, \oc8051_xiommu1/aes_top_i/reduce_nor_287/n3 ) ;   // aes_top.v(265)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_299/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(266)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_299/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_299/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_299/n2 ) ;   // aes_top.v(266)
    not (_cvpt_882, \oc8051_xiommu1/aes_top_i/reduce_nor_299/n3 ) ;   // aes_top.v(266)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_310/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(267)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_310/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_310/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_310/n2 ) ;   // aes_top.v(267)
    not (_cvpt_874, \oc8051_xiommu1/aes_top_i/reduce_nor_310/n3 ) ;   // aes_top.v(267)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_322/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(268)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_322/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_322/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_322/n2 ) ;   // aes_top.v(268)
    not (_cvpt_866, \oc8051_xiommu1/aes_top_i/reduce_nor_322/n3 ) ;   // aes_top.v(268)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_334/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(269)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_334/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_334/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_334/n2 ) ;   // aes_top.v(269)
    not (_cvpt_858, \oc8051_xiommu1/aes_top_i/reduce_nor_334/n3 ) ;   // aes_top.v(269)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_347/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/byte_counter [3]) ;   // aes_top.v(270)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_347/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_347/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_347/n2 ) ;   // aes_top.v(270)
    not (_cvpt_850, \oc8051_xiommu1/aes_top_i/reduce_nor_347/n3 ) ;   // aes_top.v(270)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_358/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(271)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_358/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_358/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_358/n2 ) ;   // aes_top.v(271)
    not (_cvpt_842, \oc8051_xiommu1/aes_top_i/reduce_nor_358/n3 ) ;   // aes_top.v(271)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_370/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(272)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_370/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_370/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_370/n2 ) ;   // aes_top.v(272)
    not (_cvpt_834, \oc8051_xiommu1/aes_top_i/reduce_nor_370/n3 ) ;   // aes_top.v(272)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_382/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(273)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_382/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_382/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_382/n2 ) ;   // aes_top.v(273)
    not (_cvpt_826, \oc8051_xiommu1/aes_top_i/reduce_nor_382/n3 ) ;   // aes_top.v(273)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_395/n2 , \oc8051_xiommu1/aes_top_i/byte_counter [2], 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(274)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_395/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_395/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_395/n2 ) ;   // aes_top.v(274)
    not (_cvpt_818, \oc8051_xiommu1/aes_top_i/reduce_nor_395/n3 ) ;   // aes_top.v(274)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_407/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(275)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_407/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_407/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_407/n2 ) ;   // aes_top.v(275)
    not (_cvpt_810, \oc8051_xiommu1/aes_top_i/reduce_nor_407/n3 ) ;   // aes_top.v(275)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_420/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(276)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_420/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_420/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_420/n2 ) ;   // aes_top.v(276)
    not (_cvpt_802, \oc8051_xiommu1/aes_top_i/reduce_nor_420/n3 ) ;   // aes_top.v(276)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_433/n2 , \oc8051_xiommu1/aes_top_i/n267 , 
        \oc8051_xiommu1/aes_top_i/n268 ) ;   // aes_top.v(277)
    or (\oc8051_xiommu1/aes_top_i/reduce_nor_433/n3 , \oc8051_xiommu1/aes_top_i/reduce_nor_433/n1 , 
        \oc8051_xiommu1/aes_top_i/reduce_nor_433/n2 ) ;   // aes_top.v(277)
    not (_cvpt_794, \oc8051_xiommu1/aes_top_i/reduce_nor_433/n3 ) ;   // aes_top.v(277)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i2  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n2 ), 
            .a(\oc8051_xiommu1/aes_ctr [1]), .b(\oc8051_xiommu1/aes_top_i/block_counter [1]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [1]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n4 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i3  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n4 ), 
            .a(\oc8051_xiommu1/aes_ctr [2]), .b(\oc8051_xiommu1/aes_top_i/block_counter [2]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [2]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n6 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i4  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n6 ), 
            .a(\oc8051_xiommu1/aes_ctr [3]), .b(\oc8051_xiommu1/aes_top_i/block_counter [3]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [3]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n8 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i5  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n8 ), 
            .a(\oc8051_xiommu1/aes_ctr [4]), .b(\oc8051_xiommu1/aes_top_i/block_counter [4]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [4]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n10 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i6  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n10 ), 
            .a(\oc8051_xiommu1/aes_ctr [5]), .b(\oc8051_xiommu1/aes_top_i/block_counter [5]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [5]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n12 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i7  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n12 ), 
            .a(\oc8051_xiommu1/aes_ctr [6]), .b(\oc8051_xiommu1/aes_top_i/block_counter [6]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [6]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n14 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i8  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n14 ), 
            .a(\oc8051_xiommu1/aes_ctr [7]), .b(\oc8051_xiommu1/aes_top_i/block_counter [7]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [7]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n16 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i9  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n16 ), 
            .a(\oc8051_xiommu1/aes_ctr [8]), .b(\oc8051_xiommu1/aes_top_i/block_counter [8]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [8]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n18 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i10  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n18 ), 
            .a(\oc8051_xiommu1/aes_ctr [9]), .b(\oc8051_xiommu1/aes_top_i/block_counter [9]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [9]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n20 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i11  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n20 ), 
            .a(\oc8051_xiommu1/aes_ctr [10]), .b(\oc8051_xiommu1/aes_top_i/block_counter [10]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [10]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n22 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i12  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n22 ), 
            .a(\oc8051_xiommu1/aes_ctr [11]), .b(\oc8051_xiommu1/aes_top_i/block_counter [11]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [11]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n24 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i13  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n24 ), 
            .a(\oc8051_xiommu1/aes_ctr [12]), .b(\oc8051_xiommu1/aes_top_i/block_counter [12]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [12]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n26 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i14  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n26 ), 
            .a(\oc8051_xiommu1/aes_ctr [13]), .b(\oc8051_xiommu1/aes_top_i/block_counter [13]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [13]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n28 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i15  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n28 ), 
            .a(\oc8051_xiommu1/aes_ctr [14]), .b(\oc8051_xiommu1/aes_top_i/block_counter [14]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [14]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n30 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i16  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n30 ), 
            .a(\oc8051_xiommu1/aes_ctr [15]), .b(\oc8051_xiommu1/aes_top_i/block_counter [15]), 
            .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [15]), .cout(\oc8051_xiommu1/aes_top_i/add_457/n32 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i17  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n32 ), 
            .a(\oc8051_xiommu1/aes_ctr [16]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [16]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n34 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i18  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n34 ), 
            .a(\oc8051_xiommu1/aes_ctr [17]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [17]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n36 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i19  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n36 ), 
            .a(\oc8051_xiommu1/aes_ctr [18]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [18]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n38 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i20  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n38 ), 
            .a(\oc8051_xiommu1/aes_ctr [19]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [19]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n40 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i21  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n40 ), 
            .a(\oc8051_xiommu1/aes_ctr [20]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [20]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n42 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i22  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n42 ), 
            .a(\oc8051_xiommu1/aes_ctr [21]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [21]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n44 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i23  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n44 ), 
            .a(\oc8051_xiommu1/aes_ctr [22]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [22]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n46 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i24  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n46 ), 
            .a(\oc8051_xiommu1/aes_ctr [23]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [23]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n48 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i25  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n48 ), 
            .a(\oc8051_xiommu1/aes_ctr [24]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [24]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n50 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i26  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n50 ), 
            .a(\oc8051_xiommu1/aes_ctr [25]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [25]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n52 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i27  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n52 ), 
            .a(\oc8051_xiommu1/aes_ctr [26]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [26]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n54 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i28  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n54 ), 
            .a(\oc8051_xiommu1/aes_ctr [27]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [27]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n56 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i29  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n56 ), 
            .a(\oc8051_xiommu1/aes_ctr [28]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [28]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n58 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i30  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n58 ), 
            .a(\oc8051_xiommu1/aes_ctr [29]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [29]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n60 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i31  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n60 ), 
            .a(\oc8051_xiommu1/aes_ctr [30]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [30]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n62 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i32  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n62 ), 
            .a(\oc8051_xiommu1/aes_ctr [31]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [31]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n64 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i33  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n64 ), 
            .a(\oc8051_xiommu1/aes_ctr [32]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [32]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n66 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i34  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n66 ), 
            .a(\oc8051_xiommu1/aes_ctr [33]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [33]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n68 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i35  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n68 ), 
            .a(\oc8051_xiommu1/aes_ctr [34]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [34]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n70 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i36  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n70 ), 
            .a(\oc8051_xiommu1/aes_ctr [35]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [35]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n72 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i37  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n72 ), 
            .a(\oc8051_xiommu1/aes_ctr [36]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [36]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n74 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i38  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n74 ), 
            .a(\oc8051_xiommu1/aes_ctr [37]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [37]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n76 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i39  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n76 ), 
            .a(\oc8051_xiommu1/aes_ctr [38]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [38]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n78 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i40  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n78 ), 
            .a(\oc8051_xiommu1/aes_ctr [39]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [39]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n80 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i41  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n80 ), 
            .a(\oc8051_xiommu1/aes_ctr [40]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [40]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n82 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i42  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n82 ), 
            .a(\oc8051_xiommu1/aes_ctr [41]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [41]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n84 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i43  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n84 ), 
            .a(\oc8051_xiommu1/aes_ctr [42]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [42]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n86 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i44  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n86 ), 
            .a(\oc8051_xiommu1/aes_ctr [43]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [43]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n88 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i45  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n88 ), 
            .a(\oc8051_xiommu1/aes_ctr [44]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [44]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n90 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i46  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n90 ), 
            .a(\oc8051_xiommu1/aes_ctr [45]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [45]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n92 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i47  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n92 ), 
            .a(\oc8051_xiommu1/aes_ctr [46]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [46]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n94 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i48  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n94 ), 
            .a(\oc8051_xiommu1/aes_ctr [47]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [47]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n96 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i49  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n96 ), 
            .a(\oc8051_xiommu1/aes_ctr [48]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [48]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n98 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i50  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n98 ), 
            .a(\oc8051_xiommu1/aes_ctr [49]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [49]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n100 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i51  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n100 ), 
            .a(\oc8051_xiommu1/aes_ctr [50]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [50]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n102 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i52  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n102 ), 
            .a(\oc8051_xiommu1/aes_ctr [51]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [51]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n104 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i53  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n104 ), 
            .a(\oc8051_xiommu1/aes_ctr [52]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [52]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n106 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i54  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n106 ), 
            .a(\oc8051_xiommu1/aes_ctr [53]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [53]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n108 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i55  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n108 ), 
            .a(\oc8051_xiommu1/aes_ctr [54]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [54]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n110 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i56  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n110 ), 
            .a(\oc8051_xiommu1/aes_ctr [55]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [55]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n112 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i57  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n112 ), 
            .a(\oc8051_xiommu1/aes_ctr [56]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [56]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n114 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i58  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n114 ), 
            .a(\oc8051_xiommu1/aes_ctr [57]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [57]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n116 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i59  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n116 ), 
            .a(\oc8051_xiommu1/aes_ctr [58]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [58]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n118 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i60  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n118 ), 
            .a(\oc8051_xiommu1/aes_ctr [59]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [59]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n120 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i61  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n120 ), 
            .a(\oc8051_xiommu1/aes_ctr [60]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [60]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n122 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i62  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n122 ), 
            .a(\oc8051_xiommu1/aes_ctr [61]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [61]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n124 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i63  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n124 ), 
            .a(\oc8051_xiommu1/aes_ctr [62]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [62]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n126 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i64  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n126 ), 
            .a(\oc8051_xiommu1/aes_ctr [63]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [63]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n128 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i65  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n128 ), 
            .a(\oc8051_xiommu1/aes_ctr [64]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [64]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n130 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i66  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n130 ), 
            .a(\oc8051_xiommu1/aes_ctr [65]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [65]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n132 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i67  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n132 ), 
            .a(\oc8051_xiommu1/aes_ctr [66]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [66]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n134 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i68  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n134 ), 
            .a(\oc8051_xiommu1/aes_ctr [67]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [67]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n136 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i69  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n136 ), 
            .a(\oc8051_xiommu1/aes_ctr [68]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [68]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n138 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i70  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n138 ), 
            .a(\oc8051_xiommu1/aes_ctr [69]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [69]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n140 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i71  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n140 ), 
            .a(\oc8051_xiommu1/aes_ctr [70]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [70]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n142 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i72  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n142 ), 
            .a(\oc8051_xiommu1/aes_ctr [71]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [71]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n144 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i73  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n144 ), 
            .a(\oc8051_xiommu1/aes_ctr [72]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [72]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n146 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i74  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n146 ), 
            .a(\oc8051_xiommu1/aes_ctr [73]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [73]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n148 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i75  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n148 ), 
            .a(\oc8051_xiommu1/aes_ctr [74]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [74]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n150 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i76  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n150 ), 
            .a(\oc8051_xiommu1/aes_ctr [75]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [75]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n152 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i77  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n152 ), 
            .a(\oc8051_xiommu1/aes_ctr [76]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [76]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n154 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i78  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n154 ), 
            .a(\oc8051_xiommu1/aes_ctr [77]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [77]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n156 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i79  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n156 ), 
            .a(\oc8051_xiommu1/aes_ctr [78]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [78]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n158 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i80  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n158 ), 
            .a(\oc8051_xiommu1/aes_ctr [79]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [79]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n160 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i81  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n160 ), 
            .a(\oc8051_xiommu1/aes_ctr [80]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [80]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n162 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i82  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n162 ), 
            .a(\oc8051_xiommu1/aes_ctr [81]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [81]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n164 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i83  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n164 ), 
            .a(\oc8051_xiommu1/aes_ctr [82]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [82]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n166 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i84  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n166 ), 
            .a(\oc8051_xiommu1/aes_ctr [83]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [83]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n168 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i85  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n168 ), 
            .a(\oc8051_xiommu1/aes_ctr [84]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [84]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n170 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i86  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n170 ), 
            .a(\oc8051_xiommu1/aes_ctr [85]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [85]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n172 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i87  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n172 ), 
            .a(\oc8051_xiommu1/aes_ctr [86]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [86]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n174 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i88  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n174 ), 
            .a(\oc8051_xiommu1/aes_ctr [87]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [87]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n176 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i89  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n176 ), 
            .a(\oc8051_xiommu1/aes_ctr [88]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [88]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n178 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i90  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n178 ), 
            .a(\oc8051_xiommu1/aes_ctr [89]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [89]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n180 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i91  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n180 ), 
            .a(\oc8051_xiommu1/aes_ctr [90]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [90]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n182 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i92  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n182 ), 
            .a(\oc8051_xiommu1/aes_ctr [91]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [91]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n184 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i93  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n184 ), 
            .a(\oc8051_xiommu1/aes_ctr [92]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [92]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n186 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i94  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n186 ), 
            .a(\oc8051_xiommu1/aes_ctr [93]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [93]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n188 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i95  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n188 ), 
            .a(\oc8051_xiommu1/aes_ctr [94]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [94]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n190 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i96  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n190 ), 
            .a(\oc8051_xiommu1/aes_ctr [95]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [95]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n192 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i97  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n192 ), 
            .a(\oc8051_xiommu1/aes_ctr [96]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [96]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n194 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i98  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n194 ), 
            .a(\oc8051_xiommu1/aes_ctr [97]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [97]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n196 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i99  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n196 ), 
            .a(\oc8051_xiommu1/aes_ctr [98]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [98]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n198 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i100  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n198 ), 
            .a(\oc8051_xiommu1/aes_ctr [99]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [99]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n200 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i101  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n200 ), 
            .a(\oc8051_xiommu1/aes_ctr [100]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [100]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n202 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i102  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n202 ), 
            .a(\oc8051_xiommu1/aes_ctr [101]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [101]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n204 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i103  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n204 ), 
            .a(\oc8051_xiommu1/aes_ctr [102]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [102]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n206 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i104  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n206 ), 
            .a(\oc8051_xiommu1/aes_ctr [103]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [103]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n208 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i105  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n208 ), 
            .a(\oc8051_xiommu1/aes_ctr [104]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [104]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n210 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i106  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n210 ), 
            .a(\oc8051_xiommu1/aes_ctr [105]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [105]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n212 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i107  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n212 ), 
            .a(\oc8051_xiommu1/aes_ctr [106]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [106]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n214 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i108  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n214 ), 
            .a(\oc8051_xiommu1/aes_ctr [107]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [107]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n216 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i109  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n216 ), 
            .a(\oc8051_xiommu1/aes_ctr [108]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [108]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n218 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i110  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n218 ), 
            .a(\oc8051_xiommu1/aes_ctr [109]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [109]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n220 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i111  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n220 ), 
            .a(\oc8051_xiommu1/aes_ctr [110]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [110]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n222 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i112  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n222 ), 
            .a(\oc8051_xiommu1/aes_ctr [111]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [111]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n224 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i113  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n224 ), 
            .a(\oc8051_xiommu1/aes_ctr [112]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [112]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n226 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i114  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n226 ), 
            .a(\oc8051_xiommu1/aes_ctr [113]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [113]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n228 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i115  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n228 ), 
            .a(\oc8051_xiommu1/aes_ctr [114]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [114]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n230 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i116  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n230 ), 
            .a(\oc8051_xiommu1/aes_ctr [115]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [115]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n232 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i117  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n232 ), 
            .a(\oc8051_xiommu1/aes_ctr [116]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [116]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n234 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i118  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n234 ), 
            .a(\oc8051_xiommu1/aes_ctr [117]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [117]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n236 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i119  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n236 ), 
            .a(\oc8051_xiommu1/aes_ctr [118]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [118]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n238 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i120  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n238 ), 
            .a(\oc8051_xiommu1/aes_ctr [119]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [119]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n240 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i121  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n240 ), 
            .a(\oc8051_xiommu1/aes_ctr [120]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [120]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n242 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i122  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n242 ), 
            .a(\oc8051_xiommu1/aes_ctr [121]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [121]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n244 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i123  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n244 ), 
            .a(\oc8051_xiommu1/aes_ctr [122]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [122]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n246 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i124  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n246 ), 
            .a(\oc8051_xiommu1/aes_ctr [123]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [123]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n248 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i125  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n248 ), 
            .a(\oc8051_xiommu1/aes_ctr [124]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [124]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n250 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i126  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n250 ), 
            .a(\oc8051_xiommu1/aes_ctr [125]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [125]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n252 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i127  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n252 ), 
            .a(\oc8051_xiommu1/aes_ctr [126]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [126]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/n254 ));   // aes_top.v(281)
    VERIFIC_FADD \oc8051_xiommu1/aes_top_i/add_457/i128  (.cin(\oc8051_xiommu1/aes_top_i/add_457/n254 ), 
            .a(\oc8051_xiommu1/aes_ctr [127]), .b(1'b0), .o(\oc8051_xiommu1/aes_top_i/aes_ctr_v [127]), 
            .cout(\oc8051_xiommu1/aes_top_i/add_457/cout ));   // aes_top.v(281)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n2 , \oc8051_xiommu1/selected_port [0], 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n1 ) ;   // oc8051_memarbiter.v(126)
    not (_cvpt_1255, \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_3/n2 ) ;   // oc8051_memarbiter.v(126)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n2 , \oc8051_xiommu1/oc8051_memarbiter_i/n5 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n1 ) ;   // oc8051_memarbiter.v(127)
    not (_cvpt_1254, \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_5/n2 ) ;   // oc8051_memarbiter.v(127)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n2 , \oc8051_xiommu1/selected_port [0], 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n1 ) ;   // oc8051_memarbiter.v(128)
    not (_cvpt_1253, \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_7/n2 ) ;   // oc8051_memarbiter.v(128)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n2 , \oc8051_xiommu1/oc8051_memarbiter_i/n5 , 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n1 ) ;   // oc8051_memarbiter.v(129)
    not (_cvpt_1252, \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_10/n2 ) ;   // oc8051_memarbiter.v(129)
    or (\oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n2 , \oc8051_xiommu1/selected_port [0], 
        \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n1 ) ;   // oc8051_memarbiter.v(150)
    not (_cvpt_1360, \oc8051_xiommu1/oc8051_memarbiter_i/reduce_nor_152/n2 ) ;   // oc8051_memarbiter.v(150)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n2  = _cvpt_3401 ? _cvpt_1411 : 1'b1;   // oc8051_page_table.v(65)
    xor (_cvpt_3402, 1'b0, _cvpt_3958) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n4  = _cvpt_3402 ? _cvpt_3958 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n2 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3403, 1'b0, _cvpt_3962) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n6  = _cvpt_3403 ? _cvpt_3962 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n4 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3404, 1'b0, _cvpt_3970) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n8  = _cvpt_3404 ? _cvpt_3970 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n6 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3405, 1'b0, _cvpt_3986) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n10  = _cvpt_3405 ? _cvpt_3986 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n8 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3406, 1'b0, \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n12  = _cvpt_3406 ? \oc8051_xiommu1/addr_out [5] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n10 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3407, 1'b0, \oc8051_xiommu1/addr_out [6]) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n14  = _cvpt_3407 ? \oc8051_xiommu1/addr_out [6] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n12 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3408, 1'b1, \oc8051_xiommu1/addr_out [7]) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n16  = _cvpt_3408 ? \oc8051_xiommu1/addr_out [7] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n14 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3409, 1'b1, _cvpt_1401) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n18  = _cvpt_3409 ? _cvpt_1401 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n16 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3410, 1'b1, _cvpt_3706) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n20  = _cvpt_3410 ? _cvpt_3706 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n18 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3411, 1'b1, _cvpt_3710) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n22  = _cvpt_3411 ? _cvpt_3710 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n20 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3412, 1'b1, _cvpt_1377) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n24  = _cvpt_3412 ? _cvpt_1377 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n22 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3413, 1'b1, _cvpt_3466) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n26  = _cvpt_3413 ? _cvpt_3466 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n24 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3414, 1'b1, _cvpt_3470) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n28  = _cvpt_3414 ? _cvpt_3470 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n26 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3415, 1'b1, _cvpt_3478) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n30  = _cvpt_3415 ? _cvpt_3478 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n28 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3416, 1'b1, _cvpt_3494) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/n4  = _cvpt_3416 ? _cvpt_3494 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_3/n30 ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n2  = _cvpt_3417 ? 1'b1 : 1'b1;   // oc8051_page_table.v(65)
    xor (_cvpt_3418, _cvpt_3958, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n4  = _cvpt_3418 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n2 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3419, _cvpt_3962, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n6  = _cvpt_3419 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n4 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3420, _cvpt_3970, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n8  = _cvpt_3420 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n6 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3421, _cvpt_3986, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n10  = _cvpt_3421 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n8 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3422, \oc8051_xiommu1/addr_out [5], 1'b0) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n12  = _cvpt_3422 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n10 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3423, \oc8051_xiommu1/addr_out [6], 1'b0) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n14  = _cvpt_3423 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n12 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3424, \oc8051_xiommu1/addr_out [7], 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n16  = _cvpt_3424 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n14 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3425, _cvpt_1401, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n18  = _cvpt_3425 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n16 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3426, _cvpt_3706, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n20  = _cvpt_3426 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n18 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3427, _cvpt_3710, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n22  = _cvpt_3427 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n20 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3428, _cvpt_1377, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n24  = _cvpt_3428 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n22 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3429, _cvpt_3466, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n26  = _cvpt_3429 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n24 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3430, _cvpt_3470, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n28  = _cvpt_3430 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n26 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3431, _cvpt_3478, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n30  = _cvpt_3431 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n28 ;   // oc8051_page_table.v(65)
    xor (_cvpt_3432, _cvpt_3494, 1'b1) ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/n5  = _cvpt_3432 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_4/n30 ;   // oc8051_page_table.v(65)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n2  = _cvpt_3433 ? _cvpt_1411 : 1'b1;   // oc8051_page_table.v(66)
    xor (_cvpt_3434, 1'b0, _cvpt_3958) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n4  = _cvpt_3434 ? _cvpt_3958 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n2 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3435, 1'b0, _cvpt_3962) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n6  = _cvpt_3435 ? _cvpt_3962 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n4 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3436, 1'b0, _cvpt_3970) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n8  = _cvpt_3436 ? _cvpt_3970 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n6 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3437, 1'b0, _cvpt_3986) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n10  = _cvpt_3437 ? _cvpt_3986 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n8 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3438, 1'b1, \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n12  = _cvpt_3438 ? \oc8051_xiommu1/addr_out [5] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n10 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3439, 1'b0, \oc8051_xiommu1/addr_out [6]) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n14  = _cvpt_3439 ? \oc8051_xiommu1/addr_out [6] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n12 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3440, 1'b1, \oc8051_xiommu1/addr_out [7]) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n16  = _cvpt_3440 ? \oc8051_xiommu1/addr_out [7] : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n14 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3441, 1'b1, _cvpt_1401) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n18  = _cvpt_3441 ? _cvpt_1401 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n16 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3442, 1'b1, _cvpt_3706) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n20  = _cvpt_3442 ? _cvpt_3706 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n18 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3443, 1'b1, _cvpt_3710) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n22  = _cvpt_3443 ? _cvpt_3710 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n20 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3444, 1'b1, _cvpt_1377) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n24  = _cvpt_3444 ? _cvpt_1377 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n22 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3445, 1'b1, _cvpt_3466) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n26  = _cvpt_3445 ? _cvpt_3466 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n24 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3446, 1'b1, _cvpt_3470) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n28  = _cvpt_3446 ? _cvpt_3470 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n26 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3447, 1'b1, _cvpt_3478) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n30  = _cvpt_3447 ? _cvpt_3478 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n28 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3448, 1'b1, _cvpt_3494) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/n7  = _cvpt_3448 ? _cvpt_3494 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_6/n30 ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n2  = _cvpt_3449 ? 1'b1 : 1'b1;   // oc8051_page_table.v(66)
    xor (_cvpt_3450, _cvpt_3958, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n4  = _cvpt_3450 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n2 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3451, _cvpt_3962, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n6  = _cvpt_3451 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n4 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3452, _cvpt_3970, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n8  = _cvpt_3452 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n6 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3453, _cvpt_3986, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n10  = _cvpt_3453 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n8 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3454, \oc8051_xiommu1/addr_out [5], 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n12  = _cvpt_3454 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n10 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3455, \oc8051_xiommu1/addr_out [6], 1'b0) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n14  = _cvpt_3455 ? 1'b0 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n12 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3456, \oc8051_xiommu1/addr_out [7], 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n16  = _cvpt_3456 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n14 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3457, _cvpt_1401, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n18  = _cvpt_3457 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n16 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3458, _cvpt_3706, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n20  = _cvpt_3458 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n18 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3459, _cvpt_3710, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n22  = _cvpt_3459 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n20 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3460, _cvpt_1377, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n24  = _cvpt_3460 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n22 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3461, _cvpt_3466, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n26  = _cvpt_3461 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n24 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3462, _cvpt_3470, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n28  = _cvpt_3462 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n26 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3463, _cvpt_3478, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n30  = _cvpt_3463 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n28 ;   // oc8051_page_table.v(66)
    xor (_cvpt_3464, _cvpt_3494, 1'b1) ;   // oc8051_page_table.v(66)
    assign \oc8051_xiommu1/oc8051_page_table_i/n8  = _cvpt_3464 ? 1'b1 : \oc8051_xiommu1/oc8051_page_table_i/LessThan_7/n30 ;   // oc8051_page_table.v(66)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n2 , _cvpt_3962, 
        _cvpt_3970) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n2 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n5 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n6 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n9 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n12 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n13 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n14 ) ;   // oc8051_page_table.v(70)
    not (_cvpt_3288, \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_20/n15 ) ;   // oc8051_page_table.v(70)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n2 , _cvpt_3962, 
        _cvpt_3970) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n2 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n5 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n6 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n9 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n12 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n13 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n14 ) ;   // oc8051_page_table.v(71)
    not (_cvpt_3272, \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_32/n15 ) ;   // oc8051_page_table.v(71)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n2 , _cvpt_3962, 
        _cvpt_3970) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n2 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n5 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n6 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n9 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n12 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n13 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n14 ) ;   // oc8051_page_table.v(72)
    not (_cvpt_3280, \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_44/n15 ) ;   // oc8051_page_table.v(72)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n2 , _cvpt_3962, 
        _cvpt_3970) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n2 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n5 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n6 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n9 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n12 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n13 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n14 ) ;   // oc8051_page_table.v(73)
    not (_cvpt_3264, \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_57/n15 ) ;   // oc8051_page_table.v(73)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n2 , \oc8051_xiommu1/oc8051_page_table_i/n59 , 
        _cvpt_3970) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n2 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n5 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n6 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n9 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n12 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n13 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n14 ) ;   // oc8051_page_table.v(74)
    not (\oc8051_xiommu1/oc8051_page_table_i/ia_pc_hi , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_69/n15 ) ;   // oc8051_page_table.v(74)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n2 , \oc8051_xiommu1/oc8051_page_table_i/n59 , 
        _cvpt_3970) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n3 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n1 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n2 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n4 , _cvpt_3986, 
        \oc8051_xiommu1/addr_out [5]) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n5 , \oc8051_xiommu1/oc8051_page_table_i/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/n12 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n6 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n4 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n5 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n7 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n3 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n6 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n8 , \oc8051_xiommu1/oc8051_page_table_i/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/n14 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n9 , \oc8051_xiommu1/oc8051_page_table_i/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/n16 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n10 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n9 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n11 , \oc8051_xiommu1/oc8051_page_table_i/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/n18 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n12 , \oc8051_xiommu1/oc8051_page_table_i/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/n20 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n13 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n12 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n14 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n13 ) ;   // oc8051_page_table.v(75)
    or (\oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n15 , \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n7 , 
        \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n14 ) ;   // oc8051_page_table.v(75)
    not (_cvpt_3256, \oc8051_xiommu1/oc8051_page_table_i/reduce_nor_82/n15 ) ;   // oc8051_page_table.v(75)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [7];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n109  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_108/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [6];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n110  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_109/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [5];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n111  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_110/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [4];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n112  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_111/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [3];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n113  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_112/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [2];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n114  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_113/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [1];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n115  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_114/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n8 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n11 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n10 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n7 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n16 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n19 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n18 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n23 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [0];   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n26 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n25 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n22 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/n116  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_115/n15 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n2  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n113  : \oc8051_xiommu1/oc8051_page_table_i/n114 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n3  = _cvpt_3706 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n1 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n4  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n111  : \oc8051_xiommu1/oc8051_page_table_i/n112 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n5  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n109  : \oc8051_xiommu1/oc8051_page_table_i/n110 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n6  = _cvpt_3706 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n4 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/wr_en  = _cvpt_3710 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_116/n3 ;   // oc8051_page_table.v(87)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n118  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_117/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n119  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_118/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n120  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_119/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n121  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_120/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n122  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_121/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n123  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_122/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n124  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_123/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n2  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n3  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n4  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n5  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n6  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n7  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n8  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n9  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n10  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n8 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n11  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n12  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n13  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n11 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n14  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n10 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n15  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n7 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n16  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n17  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n18  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n16 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n19  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n20  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n21  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n19 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n22  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n18 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n23  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n24  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n25  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n23 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n26  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n27  = _cvpt_1377 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0];   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n28  = _cvpt_3466 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n26 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n29  = _cvpt_3470 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n25 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n30  = _cvpt_3478 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n22 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/n125  = _cvpt_3494 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_124/n15 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n2  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n122  : \oc8051_xiommu1/oc8051_page_table_i/n123 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n3  = _cvpt_3706 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n1 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n4  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n120  : \oc8051_xiommu1/oc8051_page_table_i/n121 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n5  = _cvpt_1401 ? \oc8051_xiommu1/oc8051_page_table_i/n118  : \oc8051_xiommu1/oc8051_page_table_i/n119 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n6  = _cvpt_3706 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n4 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/rd_en  = _cvpt_3710 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_125/n3 ;   // oc8051_page_table.v(88)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [7] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [7];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n128  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_127/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [6] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [6];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n129  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_128/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [5] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [5];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n130  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_129/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [4] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [4];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n131  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_130/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [3] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [3];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n132  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_131/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [2] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [2];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n133  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_132/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [1] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [1];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n134  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_133/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[3] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[2] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n1 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[5] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[4] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[7] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[6] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n4 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n3 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[9] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[8] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[11] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[10] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n8 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[13] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[12] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[15] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[14] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n11 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n10 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n7 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[17] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[16] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[19] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[18] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n16 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[21] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[20] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[23] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[22] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n19 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n18 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[25] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[24] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[27] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[26] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n23 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[29] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[28] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[31] [0] : \oc8051_xiommu1/oc8051_page_table_i/wr_enabled[30] [0];   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n26 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n25 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n22 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/n135  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_134/n15 ;   // oc8051_page_table.v(92)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [7] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [7];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n144  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_143/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [6] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [6];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n145  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_144/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [5] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [5];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n146  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_145/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [4] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [4];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n147  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_146/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [3] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [3];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n148  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_147/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [2] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [2];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n149  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_148/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [1] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [1];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n150  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_149/n15 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n2  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[3] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[2] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n3  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n2  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n1 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n4  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[5] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[4] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n5  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[7] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[6] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n6  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n5  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n4 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n7  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n6  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n3 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n8  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[9] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[8] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n9  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[11] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[10] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n10  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n9  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n8 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n11  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[13] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[12] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n12  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[15] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[14] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n13  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n12  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n11 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n14  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n13  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n10 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n15  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n14  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n7 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n16  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[17] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[16] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n17  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[19] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[18] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n18  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n17  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n16 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n19  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[21] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[20] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n20  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[23] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[22] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n21  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n20  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n19 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n22  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n21  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n18 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n23  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[25] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[24] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n24  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[27] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[26] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n25  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n24  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n23 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n26  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[29] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[28] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n27  = _cvpt_1411 ? \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[31] [0] : \oc8051_xiommu1/oc8051_page_table_i/rd_enabled[30] [0];   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n28  = _cvpt_3958 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n27  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n26 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n29  = _cvpt_3962 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n28  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n25 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n30  = _cvpt_3970 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n29  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n22 ;   // oc8051_page_table.v(93)
    assign \oc8051_xiommu1/oc8051_page_table_i/n151  = _cvpt_3986 ? \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n30  : \oc8051_xiommu1/oc8051_page_table_i/Mux_150/n15 ;   // oc8051_page_table.v(93)
    not (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n3 , _cvpt_3958) ;   // oc8051_page_table.v(107)
    not (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 , _cvpt_3962) ;   // oc8051_page_table.v(107)
    not (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 , _cvpt_3970) ;   // oc8051_page_table.v(107)
    not (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 , _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n9 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n8 , 
        _cvpt_3958) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n10 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n8 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n3 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n11 , _cvpt_1411, 
        _cvpt_3958) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n12 , _cvpt_1411, 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n3 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n13 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n10 , 
        _cvpt_3962) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n14 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n10 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n15 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n12 , 
        _cvpt_3962) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n16 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n12 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n17 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n9 , 
        _cvpt_3962) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n18 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n9 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n19 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n11 , 
        _cvpt_3962) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n20 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n11 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n4 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n21 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n14 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n22 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n14 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n23 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n16 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n24 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n16 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n25 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n18 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n26 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n18 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n27 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n20 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n28 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n20 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n29 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n13 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n30 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n13 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n31 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n15 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n32 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n15 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n33 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n17 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n34 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n17 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n35 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n19 , 
        _cvpt_3970) ;   // oc8051_page_table.v(107)
    and (\oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n36 , \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n19 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n5 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1563, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n22 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1691, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n22 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1555, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n24 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1683, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n24 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1547, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n26 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1675, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n26 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1539, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n28 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1667, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n28 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1531, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n30 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1659, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n30 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1523, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n32 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1651, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n32 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1515, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n34 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1643, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n34 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1507, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n36 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1635, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n36 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1499, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n21 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1627, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n21 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1491, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n23 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1619, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n23 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1483, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n25 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1611, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n25 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1475, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n27 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1603, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n27 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1467, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n29 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1595, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n29 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1459, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n31 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1587, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n31 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1451, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n33 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1579, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n33 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    and (_cvpt_1443, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n35 , 
        _cvpt_3986) ;   // oc8051_page_table.v(107)
    and (_cvpt_1571, \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n35 , 
        \oc8051_xiommu1/oc8051_page_table_i/Decoder_161/n6 ) ;   // oc8051_page_table.v(107)
    or (_cvpt_3236, \oc8051_xiommu1/selected_port [0], \oc8051_xiommu1/oc8051_page_table_i/reduce_or_2475/n1 ) ;   // oc8051_page_table.v(129)
    
endmodule

//
// Verific Verilog Description of module oc8051_cxrom
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_symbolic_cxrom
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_ram_top
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_alu
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module termination_fsm
//

module termination_fsm (clk, rst, pout, finished);   // oc8051_tb.v(407)
    input clk;   // oc8051_tb.v(408)
    input rst;   // oc8051_tb.v(409)
    input [7:0]pout;   // oc8051_tb.v(410)
    output finished;   // oc8051_tb.v(411)
    
    wire [1:0]state;   // oc8051_tb.v(413)
    wire [1:0]state_init_next;   // oc8051_tb.v(421)
    wire [1:0]state_de_next;   // oc8051_tb.v(422)
    wire [1:0]state_ad_next;   // oc8051_tb.v(424)
    
    wire n4, n5, n7, n8, n9, n10, n11, n12, n21, n24, n26, 
        n34, n38, n39, n40, n41;
    
    not (n4, state[0]) ;   // oc8051_tb.v(419)
    not (n5, state[1]) ;   // oc8051_tb.v(419)
    nor (finished, n5, n4) ;   // oc8051_tb.v(419)
    not (n7, pout[1]) ;   // oc8051_tb.v(421)
    not (n8, pout[2]) ;   // oc8051_tb.v(421)
    not (n9, pout[3]) ;   // oc8051_tb.v(421)
    not (n10, pout[4]) ;   // oc8051_tb.v(421)
    not (n11, pout[6]) ;   // oc8051_tb.v(421)
    not (n12, pout[7]) ;   // oc8051_tb.v(421)
    nor (state_init_next[0], n12, n11, pout[5], n10, n9, n8, n7, 
        pout[0]) ;   // oc8051_tb.v(421)
    not (n21, pout[0]) ;   // oc8051_tb.v(423)
    not (n24, pout[5]) ;   // oc8051_tb.v(423)
    nor (n26, n12, pout[6], n24, pout[4], n9, n8, pout[1], n21) ;   // oc8051_tb.v(423)
    assign state_de_next[1] = state_init_next[0] ? 1'b0 : n26;   // oc8051_tb.v(423)
    nor (n34, pout[7], pout[6], pout[5], pout[4], pout[3], pout[2], 
        pout[1], pout[0]) ;   // oc8051_tb.v(425)
    assign state_ad_next[1] = n26 ? 1'b1 : n34;   // oc8051_tb.v(425)
    assign state_ad_next[0] = n26 ? 1'b0 : n34;   // oc8051_tb.v(425)
    Mux_2u_4u Mux_37 (.sel({state}), .data({1'b1, state_ad_next[1], state_de_next[1], 
            1'b0}), .o(n38));   // oc8051_tb.v(440)
    Mux_2u_4u Mux_38 (.sel({state}), .data({1'b1, state_ad_next[0], state_init_next[0], 
            state_init_next[0]}), .o(n39));   // oc8051_tb.v(440)
    assign n40 = rst ? 1'b0 : n38;   // oc8051_tb.v(441)
    assign n41 = rst ? 1'b0 : n39;   // oc8051_tb.v(441)
    VERIFIC_DFFRS i43 (.d(n41), .clk(clk), .s(1'b0), .r(1'b0), .q(state[0]));   // oc8051_tb.v(442)
    VERIFIC_DFFRS i42 (.d(n40), .clk(clk), .s(1'b0), .r(1'b0), .q(state[1]));   // oc8051_tb.v(442)
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_2u_4u
//

module Mux_2u_4u (sel, data, o);
    input [1:0]sel;
    input [3:0]data;
    output o;
    
    
    wire n1, n2;
    
    assign n1 = sel[0] ? data[1] : data[0];
    assign n2 = sel[0] ? data[3] : data[2];
    assign o = sel[1] ? n2 : n1;
    
endmodule

//
// Verific Verilog Description of module oc8051_uart_test
//

module oc8051_uart_test (clk, rst, addr, wr, wr_bit, data_in, data_out, 
            bit_out, rxd, txd, ow, intr, ack, stb);   // oc8051_uart_test.v(61)
    input clk;   // oc8051_uart_test.v(78)
    input rst;   // oc8051_uart_test.v(78)
    input [7:0]addr;   // oc8051_uart_test.v(79)
    input wr;   // oc8051_uart_test.v(78)
    input wr_bit;   // oc8051_uart_test.v(78)
    input [7:0]data_in;   // oc8051_uart_test.v(79)
    output [7:0]data_out;   // oc8051_uart_test.v(82)
    output bit_out;   // oc8051_uart_test.v(81)
    input rxd;   // oc8051_uart_test.v(78)
    output txd;   // oc8051_uart_test.v(81)
    input ow;   // oc8051_uart_test.v(78)
    output intr;   // oc8051_uart_test.v(81)
    output ack;   // oc8051_uart_test.v(81)
    input stb;   // oc8051_uart_test.v(78)
    
    wire wr_r;   // oc8051_uart_test.v(87)
    wire [7:0]addr_r;   // oc8051_uart_test.v(88)
    wire [7:0]data_in_r;   // oc8051_uart_test.v(88)
    wire brate2;   // oc8051_uart_test.v(90)
    wire pres_ow;   // oc8051_uart_test.v(95)
    wire [3:0]prescaler;   // oc8051_uart_test.v(96)
    wire [7:0]scon;   // oc8051_uart_test.v(98)
    wire [7:0]pcon;   // oc8051_uart_test.v(98)
    wire [7:0]sbuf;   // oc8051_uart_test.v(98)
    
    wire n5, n26, n27, n28, n29, n31, n32, n33, n34, n35, 
        n36, n37, n38, n89, n88, n87, n44, n45, n46, n47, 
        n48, n52, n54, n55, n57, n58;
    
    assign brate2 = 1'b0;
    oc8051_uart oc8051_uart_test (.rst(rst), .clk(clk), .bit_in(data_in[0]), 
            .data_in({data_in_r}), .wr(wr_r), .wr_bit(wr_bit), .wr_addr({addr_r}), 
            .rxd(rxd), .txd(txd), .intr(intr), .t1_ow(ow), .rclk(brate2), 
            .tclk(brate2), .pres_ow(pres_ow), .brate2(brate2), .scon({scon}), 
            .pcon({pcon}), .sbuf({sbuf}));   // oc8051_uart_test.v(100)
    assign n5 = ack ? brate2 : stb;   // oc8051_uart_test.v(111)
    VERIFIC_DFFRS i8 (.d(wr), .clk(clk), .s(brate2), .r(brate2), .q(wr_r));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i9 (.d(addr[7]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[7]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i10 (.d(addr[6]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[6]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i11 (.d(addr[5]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[5]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i12 (.d(addr[4]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[4]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i13 (.d(addr[3]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[3]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i14 (.d(addr[2]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[2]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i15 (.d(addr[1]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[1]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i16 (.d(addr[0]), .clk(clk), .s(brate2), .r(brate2), 
            .q(addr_r[0]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i17 (.d(data_in[7]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[7]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i18 (.d(data_in[6]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[6]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i19 (.d(data_in[5]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[5]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i20 (.d(data_in[4]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[4]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i21 (.d(data_in[3]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[3]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i22 (.d(data_in[2]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[2]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i23 (.d(data_in[1]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[1]));   // oc8051_uart_test.v(119)
    VERIFIC_DFFRS i24 (.d(data_in[0]), .clk(clk), .s(brate2), .r(brate2), 
            .q(data_in_r[0]));   // oc8051_uart_test.v(119)
    and (n87, rst, brate2) ;   // oc8051_uart_test.v(132)
    not (n26, prescaler[0]) ;   // oc8051_uart_test.v(126)
    not (n27, prescaler[1]) ;   // oc8051_uart_test.v(126)
    not (n28, prescaler[3]) ;   // oc8051_uart_test.v(126)
    nor (n29, n28, prescaler[2], n27, n26) ;   // oc8051_uart_test.v(126)
    add_4u_4u add_29 (.cin(brate2), .a({prescaler}), .b({brate2, brate2, 
            brate2, 1'b1}), .o({n31, n32, n33, n34}));   // oc8051_uart_test.v(130)
    assign n35 = n29 ? brate2 : n31;   // oc8051_uart_test.v(132)
    assign n36 = n29 ? brate2 : n32;   // oc8051_uart_test.v(132)
    assign n37 = n29 ? brate2 : n33;   // oc8051_uart_test.v(132)
    assign n38 = n29 ? brate2 : n34;   // oc8051_uart_test.v(132)
    VERIFIC_DFFRS i36 (.d(n36), .clk(clk), .s(rst), .r(brate2), .q(prescaler[2]));   // oc8051_uart_test.v(132)
    VERIFIC_DFFRS i38 (.d(n38), .clk(clk), .s(rst), .r(brate2), .q(prescaler[0]));   // oc8051_uart_test.v(132)
    not (n44, addr[3]) ;   // oc8051_uart_test.v(140)
    not (n45, addr[4]) ;   // oc8051_uart_test.v(140)
    not (n46, addr[7]) ;   // oc8051_uart_test.v(140)
    nor (n47, n46, addr[6], addr[5], n45, n44, addr[2], addr[1], 
        addr[0]) ;   // oc8051_uart_test.v(140)
    not (n48, addr[0]) ;   // oc8051_uart_test.v(141)
    nor (n52, n46, addr[6], addr[5], n45, n44, addr[2], addr[1], 
        n48) ;   // oc8051_uart_test.v(141)
    not (n54, addr[1]) ;   // oc8051_uart_test.v(142)
    not (n55, addr[2]) ;   // oc8051_uart_test.v(142)
    nor (n57, n46, addr[6], addr[5], addr[4], addr[3], n55, n54, 
        n48) ;   // oc8051_uart_test.v(142)
    nor (n58, n47, n52, n57) ;   // oc8051_uart_test.v(144)
    Select_4 Select_54 (.sel({n47, n52, n57, n58}), .data({scon[7], 
            sbuf[7], pcon[7], brate2}), .o(data_out[7]));   // oc8051_uart_test.v(144)
    Select_4 Select_55 (.sel({n47, n52, n57, n58}), .data({scon[6], 
            sbuf[6], pcon[6], brate2}), .o(data_out[6]));   // oc8051_uart_test.v(144)
    Select_4 Select_56 (.sel({n47, n52, n57, n58}), .data({scon[5], 
            sbuf[5], pcon[5], brate2}), .o(data_out[5]));   // oc8051_uart_test.v(144)
    Select_4 Select_57 (.sel({n47, n52, n57, n58}), .data({scon[4], 
            sbuf[4], pcon[4], brate2}), .o(data_out[4]));   // oc8051_uart_test.v(144)
    Select_4 Select_58 (.sel({n47, n52, n57, n58}), .data({scon[3], 
            sbuf[3], pcon[3], brate2}), .o(data_out[3]));   // oc8051_uart_test.v(144)
    Select_4 Select_59 (.sel({n47, n52, n57, n58}), .data({scon[2], 
            sbuf[2], pcon[2], brate2}), .o(data_out[2]));   // oc8051_uart_test.v(144)
    Select_4 Select_60 (.sel({n47, n52, n57, n58}), .data({scon[1], 
            sbuf[1], pcon[1], brate2}), .o(data_out[1]));   // oc8051_uart_test.v(144)
    Select_4 Select_61 (.sel({n47, n52, n57, n58}), .data({scon[0], 
            sbuf[0], pcon[0], brate2}), .o(data_out[0]));   // oc8051_uart_test.v(144)
    Mux_3u_8u Mux_62 (.sel({addr[2:0]}), .data({scon}), .o(bit_out));   // oc8051_uart_test.v(147)
    VERIFIC_DFFRS i6 (.d(n5), .clk(clk), .s(brate2), .r(brate2), .q(ack));   // oc8051_uart_test.v(112)
    not (n88, brate2) ;   // oc8051_uart_test.v(132)
    and (n89, rst, n88) ;   // oc8051_uart_test.v(132)
    VERIFIC_DFFRS i35 (.d(n35), .clk(clk), .s(n87), .r(n89), .q(prescaler[3]));   // oc8051_uart_test.v(132)
    VERIFIC_DFFRS i37 (.d(n37), .clk(clk), .s(n87), .r(n89), .q(prescaler[1]));   // oc8051_uart_test.v(132)
    VERIFIC_DFFRS i39 (.d(n29), .clk(clk), .s(n87), .r(n89), .q(pres_ow));   // oc8051_uart_test.v(132)
    
endmodule

//
// Verific Verilog Description of module oc8051_uart
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of OPERATOR add_4u_4u
//

module add_4u_4u (cin, a, b, o, cout);
    input cin;
    input [3:0]a;
    input [3:0]b;
    output [3:0]o;
    output cout;
    
    
    wire n2, n4, n6;
    
    VERIFIC_FADD i1 (.cin(cin), .a(a[0]), .b(b[0]), .o(o[0]), .cout(n2));
    VERIFIC_FADD i2 (.cin(n2), .a(a[1]), .b(b[1]), .o(o[1]), .cout(n4));
    VERIFIC_FADD i3 (.cin(n4), .a(a[2]), .b(b[2]), .o(o[2]), .cout(n6));
    VERIFIC_FADD i4 (.cin(n6), .a(a[3]), .b(b[3]), .o(o[3]), .cout(cout));
    
endmodule

//
// Verific Verilog Description of OPERATOR Select_4
//

module Select_4 (sel, data, o);
    input [3:0]sel;
    input [3:0]data;
    output o;
    
    
    wire n1, n2, n3, n4, n5, n6;
    
    and (n1, data[0], sel[0]) ;
    and (n2, data[1], sel[1]) ;
    and (n3, data[2], sel[2]) ;
    and (n4, data[3], sel[3]) ;
    or (n5, n1, n2) ;
    or (n6, n3, n4) ;
    or (o, n5, n6) ;
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_3u_8u
//

module Mux_3u_8u (sel, data, o);
    input [2:0]sel;
    input [7:0]data;
    output o;
    
    
    wire n1, n2, n3, n4, n5, n6;
    
    assign n1 = sel[0] ? data[1] : data[0];
    assign n2 = sel[0] ? data[3] : data[2];
    assign n3 = sel[1] ? n2 : n1;
    assign n4 = sel[0] ? data[5] : data[4];
    assign n5 = sel[0] ? data[7] : data[6];
    assign n6 = sel[1] ? n5 : n4;
    assign o = sel[2] ? n6 : n3;
    
endmodule

//
// Verific Verilog Description of module oc8051_alu_src_sel
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_comp
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_rom
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_cy_select
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_indi_addr
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_memory_interface
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_sfr
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_priv_lvl
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module sha_top
//

module sha_top (clk, rst, wr, addr, data_in, data_out, ack, stb, 
            in_addr_range, xram_addr, xram_data_out, xram_data_in, xram_ack, 
            xram_stb, xram_wr, sha_state, sha_rdaddr, sha_wraddr, 
            sha_len, sha_step, sha_core_assumps_valid);   // sha_top.v(12)
    input clk;   // sha_top.v(49)
    input rst;   // sha_top.v(49)
    input wr;   // sha_top.v(49)
    input [15:0]addr;   // sha_top.v(51)
    input [7:0]data_in;   // sha_top.v(50)
    output [7:0]data_out;   // sha_top.v(52)
    output ack;   // sha_top.v(53)
    input stb;   // sha_top.v(49)
    output in_addr_range;   // sha_top.v(54)
    output [15:0]xram_addr;   // sha_top.v(56)
    output [7:0]xram_data_out;   // sha_top.v(57)
    input [7:0]xram_data_in;   // sha_top.v(58)
    input xram_ack;   // sha_top.v(59)
    output xram_stb;   // sha_top.v(60)
    output xram_wr;   // sha_top.v(61)
    output [2:0]sha_state;   // sha_top.v(63)
    output [15:0]sha_rdaddr;   // sha_top.v(64)
    output [15:0]sha_wraddr;   // sha_top.v(64)
    output [15:0]sha_len;   // sha_top.v(64)
    output sha_step;   // sha_top.v(65)
    output sha_core_assumps_valid;   // sha_top.v(66)
    
    wire sha_state_idle;   // sha_top.v(92)
    wire sha_state_read_data;   // sha_top.v(93)
    wire sha_state_op1;   // sha_top.v(94)
    wire sha_state_op2;   // sha_top.v(95)
    wire sel_reg_start;   // sha_top.v(99)
    wire sel_reg_state;   // sha_top.v(100)
    wire sel_reg_rd_addr;   // sha_top.v(101)
    wire sel_reg_wr_addr;   // sha_top.v(102)
    wire sel_reg_len;   // sha_top.v(103)
    wire wren;   // sha_top.v(104)
    wire [2:0]sha_state_next;   // sha_top.v(116)
    wire [2:0]sha_state_next_idle;   // sha_top.v(118)
    wire [2:0]sha_state_next_read_data;   // sha_top.v(119)
    wire [2:0]sha_state_next_op2;   // sha_top.v(121)
    wire [2:0]sha_state_next_write_data;   // sha_top.v(122)
    wire [5:0]byte_counter;   // sha_top.v(146)
    wire [5:0]byte_counter_next;   // sha_top.v(147)
    wire [5:0]byte_counter_next_rw;   // sha_top.v(148)
    wire [15:0]reg_bytes_read;   // sha_top.v(156)
    wire [15:0]bytes_read_next;   // sha_top.v(157)
    wire [15:0]block_counter;   // sha_top.v(163)
    wire [15:0]block_counter_next;   // sha_top.v(164)
    wire reading_last_byte;   // sha_top.v(170)
    wire sha_more_blocks;   // sha_top.v(174)
    wire sha_finished;   // sha_top.v(175)
    wire [511:0]sha_core_block_read_data_next;   // sha_top.v(178)
    wire [511:0]sha_core_block_next;   // sha_top.v(245)
    wire writing_last_byte;   // sha_top.v(250)
    wire write_last_byte_acked;   // sha_top.v(251)
    wire [7:0]data_out_rd_addr;   // sha_top.v(254)
    wire [7:0]data_out_wr_addr;   // sha_top.v(255)
    wire [7:0]data_out_len;   // sha_top.v(256)
    wire sha_core_rst_n;   // sha_top.v(312)
    wire sha_core_init;   // sha_top.v(314)
    wire sha_core_next;   // sha_top.v(316)
    wire sha_core_ready;   // sha_top.v(318)
    wire sha_core_ready_r;   // sha_top.v(320)
    wire sha_core_digest_valid;   // sha_top.v(322)
    wire [511:0]sha_core_block;   // sha_top.v(324)
    wire [159:0]sha_core_digest;   // sha_top.v(326)
    wire [159:0]sha_reg_digest;   // sha_top.v(328)
    wire [159:0]sha_reg_digest_next;   // sha_top.v(330)
    
    wire n4, n5, n9, n11, n16, n18, n19, n20, n21, n22, 
        n23, n24, n26, n35, n44, n64, n65, n67, n68, n69, 
        n70, n71, n72, n73, n74, n75, n79, n80, n81, n84, 
        n89, n90, n91, n92, n93, n94, n102, n103, n104, n105, 
        n106, n107, n108, n109, n110, n111, n112, n113, n114, 
        n115, n122, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, 
        n150, n151, n152, n153, n154, n155, n156, n174, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, 
        n187, n188, n189, n190, n191, n192, n193, n194, n195, 
        n196, n214, n215, n216, n217, n218, n219, n221, n222, 
        n223, n224, n225, n226, n227, n228, n229, n230, n231, 
        n232, n233, n234, n235, n236, n237, n240, n242, n250, 
        n264, n278, n291, n305, n318, n331, n343, n357, n370, 
        n383, n395, n408, n420, n432, n443, n457, n470, n483, 
        n495, n508, n520, n532, n543, n556, n568, n580, n591, 
        n603, n614, n625, n635, n649, n662, n675, n687, n700, 
        n712, n724, n735, n748, n760, n772, n783, n806, n817, 
        n827, n840, n852, n864, n875, n887, n898, n909, n919, 
        n931, n942, n953, n963, n974, n984, n994, n1003, n1012, 
        n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
        n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
        n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
        n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, 
        n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
        n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
        n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
        n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
        n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
        n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
        n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
        n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
        n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
        n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
        n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
        n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
        n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
        n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
        n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
        n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
        n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
        n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
        n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
        n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
        n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
        n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
        n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
        n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
        n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
        n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
        n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
        n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
        n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
        n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
        n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
        n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
        n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
        n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
        n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
        n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
        n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
        n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
        n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
        n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
        n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
        n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
        n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
        n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
        n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
        n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
        n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
        n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
        n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
        n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
        n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
        n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
        n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
        n1517, n1518, n1519, n1520, n1521, n1522, n1523, n2041, 
        n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
        n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
        n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2073, 
        n2074, n2075, n2077, n2078, n2081, n2250, n2251, n2252, 
        n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
        n2261, n2262, n2263, n2264, n2265, n2267, n2268, n2269, 
        n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
        n2278, n2279, n2280, n2281, n2282, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2376, n2377, n2378, 
        n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
        n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
        n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
        n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
        n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
        n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
        n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
        n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
        n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
        n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
        n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
        n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
        n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
        n2515, n2516, n2517, n2518, n2519, n2530, n2531, n2532, 
        n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
        n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
        n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
        n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
        n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
        n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
        n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
        n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
        n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
        n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
        n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
        n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
        n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
        n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
        n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
        n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
        n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
        n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
        n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
        n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
        n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
        n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
        n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
        n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
        n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
        n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
        n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
        n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
        n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, 
        n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
        n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
        n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
        n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
        n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, 
        n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
        n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
        n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
        n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
        n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, 
        n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
        n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
        n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
        n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
        n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
        n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
        n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
        n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
        n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
        n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
        n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, 
        n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
        n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
        n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
        n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
        n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, 
        n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
        n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
        n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
        n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
        n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
        n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
        n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
        n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
        n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
        n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
        n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
        n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, 
        n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
        n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
        n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
        n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
        n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, 
        n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
        n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
        n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
        n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
        n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
        n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
        n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
        n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
        n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
        n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
        n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
        n3237, n3238, n3239, n3240, n3241, n3242, n3243;
    
    assign sha_core_assumps_valid = 1'b1;
    LessThan_16u_16u LessThan_3 (.cin(1'b1), .a({16'b1111111000000000}), 
            .b({addr}), .o(n4));   // sha_top.v(84)
    LessThan_16u_16u LessThan_4 (.cin(1'b0), .a({addr}), .b({16'b1111111000010000}), 
            .o(n5));   // sha_top.v(84)
    and (in_addr_range, n4, n5) ;   // sha_top.v(84)
    and (ack, stb, in_addr_range) ;   // sha_top.v(85)
    nor (sha_state_idle, sha_state[2], sha_state[1], sha_state[0]) ;   // sha_top.v(92)
    not (n9, sha_state[0]) ;   // sha_top.v(93)
    nor (sha_state_read_data, sha_state[2], sha_state[1], n9) ;   // sha_top.v(93)
    not (n11, sha_state[1]) ;   // sha_top.v(94)
    nor (sha_state_op1, sha_state[2], n11, sha_state[0]) ;   // sha_top.v(94)
    nor (sha_state_op2, sha_state[2], n11, n9) ;   // sha_top.v(95)
    not (n16, sha_state[2]) ;   // sha_top.v(96)
    nor (xram_wr, n16, sha_state[1], sha_state[0]) ;   // sha_top.v(96)
    not (n18, addr[9]) ;   // sha_top.v(99)
    not (n19, addr[10]) ;   // sha_top.v(99)
    not (n20, addr[11]) ;   // sha_top.v(99)
    not (n21, addr[12]) ;   // sha_top.v(99)
    not (n22, addr[13]) ;   // sha_top.v(99)
    not (n23, addr[14]) ;   // sha_top.v(99)
    not (n24, addr[15]) ;   // sha_top.v(99)
    nor (sel_reg_start, n24, n23, n22, n21, n20, n19, n18, addr[8], 
        addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], addr[1], 
        addr[0]) ;   // sha_top.v(99)
    not (n26, addr[0]) ;   // sha_top.v(100)
    nor (sel_reg_state, n24, n23, n22, n21, n20, n19, n18, addr[8], 
        addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], addr[1], 
        n26) ;   // sha_top.v(100)
    not (n35, addr[1]) ;   // sha_top.v(101)
    nor (sel_reg_rd_addr, n24, n23, n22, n21, n20, n19, n18, 
        addr[8], addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], 
        n35) ;   // sha_top.v(101)
    not (n44, addr[2]) ;   // sha_top.v(102)
    nor (sel_reg_wr_addr, n24, n23, n22, n21, n20, n19, n18, 
        addr[8], addr[7], addr[6], addr[5], addr[4], addr[3], n44, 
        addr[1]) ;   // sha_top.v(102)
    nor (sel_reg_len, n24, n23, n22, n21, n20, n19, n18, addr[8], 
        addr[7], addr[6], addr[5], addr[4], addr[3], n44, n35) ;   // sha_top.v(103)
    and (wren, wr, sha_state_idle) ;   // sha_top.v(104)
    and (n64, sel_reg_start, data_in[0]) ;   // sha_top.v(106)
    and (n65, n64, stb) ;   // sha_top.v(106)
    and (sha_state_next_idle[0], n65, wren) ;   // sha_top.v(106)
    assign n67 = sha_state_op2 ? sha_finished : sha_state_next_write_data[2];   // sha_top.v(129)
    assign n68 = sha_state_op2 ? sha_state_next_op2[1] : 1'b0;   // sha_top.v(129)
    assign n69 = sha_state_op2 ? sha_state_next_op2[0] : 1'b0;   // sha_top.v(129)
    assign n70 = sha_state_op1 ? 1'b0 : n67;   // sha_top.v(129)
    assign n71 = sha_state_op1 ? 1'b1 : n68;   // sha_top.v(129)
    assign n72 = sha_state_op1 ? 1'b1 : n69;   // sha_top.v(129)
    assign n73 = sha_state_read_data ? 1'b0 : n70;   // sha_top.v(129)
    assign n74 = sha_state_read_data ? sha_state_next_read_data[1] : n71;   // sha_top.v(129)
    assign n75 = sha_state_read_data ? sha_state_next_read_data[0] : n72;   // sha_top.v(129)
    assign sha_state_next[2] = sha_state_idle ? 1'b0 : n73;   // sha_top.v(129)
    assign sha_state_next[1] = sha_state_idle ? 1'b0 : n74;   // sha_top.v(129)
    assign sha_state_next[0] = sha_state_idle ? sha_state_next_idle[0] : n75;   // sha_top.v(129)
    xor (n79, sha_state[0], sha_state_next[0]) ;   // sha_top.v(131)
    xor (n80, sha_state[1], sha_state_next[1]) ;   // sha_top.v(131)
    xor (n81, sha_state[2], sha_state_next[2]) ;   // sha_top.v(131)
    or (sha_step, n81, n80, n79) ;   // sha_top.v(131)
    not (sha_state_next_read_data[0], sha_state_next_read_data[1]) ;   // sha_top.v(136)
    not (n84, sha_more_blocks) ;   // sha_top.v(141)
    assign sha_state_next_op2[1] = sha_finished ? 1'b0 : n84;   // sha_top.v(141)
    not (sha_state_next_op2[0], sha_finished) ;   // sha_top.v(141)
    not (sha_state_next_write_data[2], write_last_byte_acked) ;   // sha_top.v(143)
    add_6u_6u add_87 (.cin(1'b0), .a({byte_counter}), .b({6'b000001}), 
            .o({n89, n90, n91, n92, n93, n94}));   // sha_top.v(149)
    assign byte_counter_next_rw[5] = xram_ack ? n89 : byte_counter[5];   // sha_top.v(149)
    assign byte_counter_next_rw[4] = xram_ack ? n90 : byte_counter[4];   // sha_top.v(149)
    assign byte_counter_next_rw[3] = xram_ack ? n91 : byte_counter[3];   // sha_top.v(149)
    assign byte_counter_next_rw[2] = xram_ack ? n92 : byte_counter[2];   // sha_top.v(149)
    assign byte_counter_next_rw[1] = xram_ack ? n93 : byte_counter[1];   // sha_top.v(149)
    assign byte_counter_next_rw[0] = xram_ack ? n94 : byte_counter[0];   // sha_top.v(149)
    or (n102, sha_state_idle, sha_state_op1) ;   // sha_top.v(151)
    or (n103, n102, sha_state_op2) ;   // sha_top.v(151)
    assign n104 = xram_wr ? byte_counter_next_rw[5] : byte_counter[5];   // sha_top.v(153)
    assign n105 = xram_wr ? byte_counter_next_rw[4] : byte_counter[4];   // sha_top.v(153)
    assign n106 = xram_wr ? byte_counter_next_rw[3] : byte_counter[3];   // sha_top.v(153)
    assign n107 = xram_wr ? byte_counter_next_rw[2] : byte_counter[2];   // sha_top.v(153)
    assign n108 = xram_wr ? byte_counter_next_rw[1] : byte_counter[1];   // sha_top.v(153)
    assign n109 = xram_wr ? byte_counter_next_rw[0] : byte_counter[0];   // sha_top.v(153)
    assign n110 = sha_state_read_data ? byte_counter_next_rw[5] : n104;   // sha_top.v(153)
    assign n111 = sha_state_read_data ? byte_counter_next_rw[4] : n105;   // sha_top.v(153)
    assign n112 = sha_state_read_data ? byte_counter_next_rw[3] : n106;   // sha_top.v(153)
    assign n113 = sha_state_read_data ? byte_counter_next_rw[2] : n107;   // sha_top.v(153)
    assign n114 = sha_state_read_data ? byte_counter_next_rw[1] : n108;   // sha_top.v(153)
    assign n115 = sha_state_read_data ? byte_counter_next_rw[0] : n109;   // sha_top.v(153)
    assign byte_counter_next[5] = n103 ? 1'b0 : n110;   // sha_top.v(153)
    assign byte_counter_next[4] = n103 ? 1'b0 : n111;   // sha_top.v(153)
    assign byte_counter_next[3] = n103 ? 1'b0 : n112;   // sha_top.v(153)
    assign byte_counter_next[2] = n103 ? 1'b0 : n113;   // sha_top.v(153)
    assign byte_counter_next[1] = n103 ? 1'b0 : n114;   // sha_top.v(153)
    assign byte_counter_next[0] = n103 ? 1'b0 : n115;   // sha_top.v(153)
    and (n122, sha_state_read_data, xram_ack) ;   // sha_top.v(160)
    add_16u_16u add_116 (.cin(1'b0), .a({reg_bytes_read}), .b({16'b0000000000000001}), 
            .o({n124, n125, n126, n127, n128, n129, n130, n131, 
            n132, n133, n134, n135, n136, n137, n138, n139}));   // sha_top.v(160)
    assign n141 = n122 ? n124 : reg_bytes_read[15];   // sha_top.v(160)
    assign n142 = n122 ? n125 : reg_bytes_read[14];   // sha_top.v(160)
    assign n143 = n122 ? n126 : reg_bytes_read[13];   // sha_top.v(160)
    assign n144 = n122 ? n127 : reg_bytes_read[12];   // sha_top.v(160)
    assign n145 = n122 ? n128 : reg_bytes_read[11];   // sha_top.v(160)
    assign n146 = n122 ? n129 : reg_bytes_read[10];   // sha_top.v(160)
    assign n147 = n122 ? n130 : reg_bytes_read[9];   // sha_top.v(160)
    assign n148 = n122 ? n131 : reg_bytes_read[8];   // sha_top.v(160)
    assign n149 = n122 ? n132 : reg_bytes_read[7];   // sha_top.v(160)
    assign n150 = n122 ? n133 : reg_bytes_read[6];   // sha_top.v(160)
    assign n151 = n122 ? n134 : reg_bytes_read[5];   // sha_top.v(160)
    assign n152 = n122 ? n135 : reg_bytes_read[4];   // sha_top.v(160)
    assign n153 = n122 ? n136 : reg_bytes_read[3];   // sha_top.v(160)
    assign n154 = n122 ? n137 : reg_bytes_read[2];   // sha_top.v(160)
    assign n155 = n122 ? n138 : reg_bytes_read[1];   // sha_top.v(160)
    assign n156 = n122 ? n139 : reg_bytes_read[0];   // sha_top.v(160)
    assign bytes_read_next[15] = sha_state_idle ? 1'b0 : n141;   // sha_top.v(160)
    assign bytes_read_next[14] = sha_state_idle ? 1'b0 : n142;   // sha_top.v(160)
    assign bytes_read_next[13] = sha_state_idle ? 1'b0 : n143;   // sha_top.v(160)
    assign bytes_read_next[12] = sha_state_idle ? 1'b0 : n144;   // sha_top.v(160)
    assign bytes_read_next[11] = sha_state_idle ? 1'b0 : n145;   // sha_top.v(160)
    assign bytes_read_next[10] = sha_state_idle ? 1'b0 : n146;   // sha_top.v(160)
    assign bytes_read_next[9] = sha_state_idle ? 1'b0 : n147;   // sha_top.v(160)
    assign bytes_read_next[8] = sha_state_idle ? 1'b0 : n148;   // sha_top.v(160)
    assign bytes_read_next[7] = sha_state_idle ? 1'b0 : n149;   // sha_top.v(160)
    assign bytes_read_next[6] = sha_state_idle ? 1'b0 : n150;   // sha_top.v(160)
    assign bytes_read_next[5] = sha_state_idle ? 1'b0 : n151;   // sha_top.v(160)
    assign bytes_read_next[4] = sha_state_idle ? 1'b0 : n152;   // sha_top.v(160)
    assign bytes_read_next[3] = sha_state_idle ? 1'b0 : n153;   // sha_top.v(160)
    assign bytes_read_next[2] = sha_state_idle ? 1'b0 : n154;   // sha_top.v(160)
    assign bytes_read_next[1] = sha_state_idle ? 1'b0 : n155;   // sha_top.v(160)
    assign bytes_read_next[0] = sha_state_idle ? 1'b0 : n156;   // sha_top.v(160)
    and (n174, sha_state_op2, sha_more_blocks) ;   // sha_top.v(167)
    add_10u_10u add_152 (.cin(1'b0), .a({block_counter[15:6]}), .b({10'b0000000001}), 
            .o({n176, n177, n178, n179, n180, n181, n182, n183, 
            n184, n185}));   // sha_top.v(167)
    assign n187 = n174 ? n176 : block_counter[15];   // sha_top.v(167)
    assign n188 = n174 ? n177 : block_counter[14];   // sha_top.v(167)
    assign n189 = n174 ? n178 : block_counter[13];   // sha_top.v(167)
    assign n190 = n174 ? n179 : block_counter[12];   // sha_top.v(167)
    assign n191 = n174 ? n180 : block_counter[11];   // sha_top.v(167)
    assign n192 = n174 ? n181 : block_counter[10];   // sha_top.v(167)
    assign n193 = n174 ? n182 : block_counter[9];   // sha_top.v(167)
    assign n194 = n174 ? n183 : block_counter[8];   // sha_top.v(167)
    assign n195 = n174 ? n184 : block_counter[7];   // sha_top.v(167)
    assign n196 = n174 ? n185 : block_counter[6];   // sha_top.v(167)
    assign block_counter_next[15] = sha_state_idle ? 1'b0 : n187;   // sha_top.v(167)
    assign block_counter_next[14] = sha_state_idle ? 1'b0 : n188;   // sha_top.v(167)
    assign block_counter_next[13] = sha_state_idle ? 1'b0 : n189;   // sha_top.v(167)
    assign block_counter_next[12] = sha_state_idle ? 1'b0 : n190;   // sha_top.v(167)
    assign block_counter_next[11] = sha_state_idle ? 1'b0 : n191;   // sha_top.v(167)
    assign block_counter_next[10] = sha_state_idle ? 1'b0 : n192;   // sha_top.v(167)
    assign block_counter_next[9] = sha_state_idle ? 1'b0 : n193;   // sha_top.v(167)
    assign block_counter_next[8] = sha_state_idle ? 1'b0 : n194;   // sha_top.v(167)
    assign block_counter_next[7] = sha_state_idle ? 1'b0 : n195;   // sha_top.v(167)
    assign block_counter_next[6] = sha_state_idle ? 1'b0 : n196;   // sha_top.v(167)
    assign block_counter_next[5] = sha_state_idle ? 1'b0 : block_counter[5];   // sha_top.v(167)
    assign block_counter_next[4] = sha_state_idle ? 1'b0 : block_counter[4];   // sha_top.v(167)
    assign block_counter_next[3] = sha_state_idle ? 1'b0 : block_counter[3];   // sha_top.v(167)
    assign block_counter_next[2] = sha_state_idle ? 1'b0 : block_counter[2];   // sha_top.v(167)
    assign block_counter_next[1] = sha_state_idle ? 1'b0 : block_counter[1];   // sha_top.v(167)
    assign block_counter_next[0] = sha_state_idle ? 1'b0 : block_counter[0];   // sha_top.v(167)
    not (n214, byte_counter[0]) ;   // sha_top.v(170)
    not (n215, byte_counter[1]) ;   // sha_top.v(170)
    not (n216, byte_counter[2]) ;   // sha_top.v(170)
    not (n217, byte_counter[3]) ;   // sha_top.v(170)
    not (n218, byte_counter[4]) ;   // sha_top.v(170)
    not (n219, byte_counter[5]) ;   // sha_top.v(170)
    nor (n250, n219, n218, n217, n216, n215, n214) ;   // sha_top.v(170)
    xor (n221, bytes_read_next[0], sha_len[0]) ;   // sha_top.v(170)
    xor (n222, bytes_read_next[1], sha_len[1]) ;   // sha_top.v(170)
    xor (n223, bytes_read_next[2], sha_len[2]) ;   // sha_top.v(170)
    xor (n224, bytes_read_next[3], sha_len[3]) ;   // sha_top.v(170)
    xor (n225, bytes_read_next[4], sha_len[4]) ;   // sha_top.v(170)
    xor (n226, bytes_read_next[5], sha_len[5]) ;   // sha_top.v(170)
    xor (n227, bytes_read_next[6], sha_len[6]) ;   // sha_top.v(170)
    xor (n228, bytes_read_next[7], sha_len[7]) ;   // sha_top.v(170)
    xor (n229, bytes_read_next[8], sha_len[8]) ;   // sha_top.v(170)
    xor (n230, bytes_read_next[9], sha_len[9]) ;   // sha_top.v(170)
    xor (n231, bytes_read_next[10], sha_len[10]) ;   // sha_top.v(170)
    xor (n232, bytes_read_next[11], sha_len[11]) ;   // sha_top.v(170)
    xor (n233, bytes_read_next[12], sha_len[12]) ;   // sha_top.v(170)
    xor (n234, bytes_read_next[13], sha_len[13]) ;   // sha_top.v(170)
    xor (n235, bytes_read_next[14], sha_len[14]) ;   // sha_top.v(170)
    xor (n236, bytes_read_next[15], sha_len[15]) ;   // sha_top.v(170)
    nor (n237, n236, n235, n234, n233, n232, n231, n230, n229, 
        n228, n227, n226, n225, n224, n223, n222, n221) ;   // sha_top.v(170)
    or (reading_last_byte, n250, n237) ;   // sha_top.v(170)
    and (sha_state_next_read_data[1], reading_last_byte, xram_ack) ;   // sha_top.v(171)
    LessThan_16u_16u LessThan_207 (.cin(1'b0), .a({reg_bytes_read}), .b({sha_len}), 
            .o(n240));   // sha_top.v(174)
    and (sha_more_blocks, sha_core_digest_valid, n240) ;   // sha_top.v(174)
    not (n242, n240) ;   // sha_top.v(175)
    and (sha_finished, sha_core_digest_valid, n242) ;   // sha_top.v(175)
    assign sha_core_block_read_data_next[7] = n250 ? xram_data_in[7] : sha_core_block[7];   // sha_top.v(180)
    assign sha_core_block_read_data_next[6] = n250 ? xram_data_in[6] : sha_core_block[6];   // sha_top.v(180)
    assign sha_core_block_read_data_next[5] = n250 ? xram_data_in[5] : sha_core_block[5];   // sha_top.v(180)
    assign sha_core_block_read_data_next[4] = n250 ? xram_data_in[4] : sha_core_block[4];   // sha_top.v(180)
    assign sha_core_block_read_data_next[3] = n250 ? xram_data_in[3] : sha_core_block[3];   // sha_top.v(180)
    assign sha_core_block_read_data_next[2] = n250 ? xram_data_in[2] : sha_core_block[2];   // sha_top.v(180)
    assign sha_core_block_read_data_next[1] = n250 ? xram_data_in[1] : sha_core_block[1];   // sha_top.v(180)
    assign sha_core_block_read_data_next[0] = n250 ? xram_data_in[0] : sha_core_block[0];   // sha_top.v(180)
    nor (n264, n219, n218, n217, n216, n215, byte_counter[0]) ;   // sha_top.v(181)
    assign sha_core_block_read_data_next[15] = n264 ? xram_data_in[7] : sha_core_block[15];   // sha_top.v(181)
    assign sha_core_block_read_data_next[14] = n264 ? xram_data_in[6] : sha_core_block[14];   // sha_top.v(181)
    assign sha_core_block_read_data_next[13] = n264 ? xram_data_in[5] : sha_core_block[13];   // sha_top.v(181)
    assign sha_core_block_read_data_next[12] = n264 ? xram_data_in[4] : sha_core_block[12];   // sha_top.v(181)
    assign sha_core_block_read_data_next[11] = n264 ? xram_data_in[3] : sha_core_block[11];   // sha_top.v(181)
    assign sha_core_block_read_data_next[10] = n264 ? xram_data_in[2] : sha_core_block[10];   // sha_top.v(181)
    assign sha_core_block_read_data_next[9] = n264 ? xram_data_in[1] : sha_core_block[9];   // sha_top.v(181)
    assign sha_core_block_read_data_next[8] = n264 ? xram_data_in[0] : sha_core_block[8];   // sha_top.v(181)
    nor (n278, n219, n218, n217, n216, byte_counter[1], n214) ;   // sha_top.v(182)
    assign sha_core_block_read_data_next[23] = n278 ? xram_data_in[7] : sha_core_block[23];   // sha_top.v(182)
    assign sha_core_block_read_data_next[22] = n278 ? xram_data_in[6] : sha_core_block[22];   // sha_top.v(182)
    assign sha_core_block_read_data_next[21] = n278 ? xram_data_in[5] : sha_core_block[21];   // sha_top.v(182)
    assign sha_core_block_read_data_next[20] = n278 ? xram_data_in[4] : sha_core_block[20];   // sha_top.v(182)
    assign sha_core_block_read_data_next[19] = n278 ? xram_data_in[3] : sha_core_block[19];   // sha_top.v(182)
    assign sha_core_block_read_data_next[18] = n278 ? xram_data_in[2] : sha_core_block[18];   // sha_top.v(182)
    assign sha_core_block_read_data_next[17] = n278 ? xram_data_in[1] : sha_core_block[17];   // sha_top.v(182)
    assign sha_core_block_read_data_next[16] = n278 ? xram_data_in[0] : sha_core_block[16];   // sha_top.v(182)
    nor (n291, n219, n218, n217, n216, byte_counter[1], byte_counter[0]) ;   // sha_top.v(183)
    assign sha_core_block_read_data_next[31] = n291 ? xram_data_in[7] : sha_core_block[31];   // sha_top.v(183)
    assign sha_core_block_read_data_next[30] = n291 ? xram_data_in[6] : sha_core_block[30];   // sha_top.v(183)
    assign sha_core_block_read_data_next[29] = n291 ? xram_data_in[5] : sha_core_block[29];   // sha_top.v(183)
    assign sha_core_block_read_data_next[28] = n291 ? xram_data_in[4] : sha_core_block[28];   // sha_top.v(183)
    assign sha_core_block_read_data_next[27] = n291 ? xram_data_in[3] : sha_core_block[27];   // sha_top.v(183)
    assign sha_core_block_read_data_next[26] = n291 ? xram_data_in[2] : sha_core_block[26];   // sha_top.v(183)
    assign sha_core_block_read_data_next[25] = n291 ? xram_data_in[1] : sha_core_block[25];   // sha_top.v(183)
    assign sha_core_block_read_data_next[24] = n291 ? xram_data_in[0] : sha_core_block[24];   // sha_top.v(183)
    nor (n305, n219, n218, n217, byte_counter[2], n215, n214) ;   // sha_top.v(184)
    assign sha_core_block_read_data_next[39] = n305 ? xram_data_in[7] : sha_core_block[39];   // sha_top.v(184)
    assign sha_core_block_read_data_next[38] = n305 ? xram_data_in[6] : sha_core_block[38];   // sha_top.v(184)
    assign sha_core_block_read_data_next[37] = n305 ? xram_data_in[5] : sha_core_block[37];   // sha_top.v(184)
    assign sha_core_block_read_data_next[36] = n305 ? xram_data_in[4] : sha_core_block[36];   // sha_top.v(184)
    assign sha_core_block_read_data_next[35] = n305 ? xram_data_in[3] : sha_core_block[35];   // sha_top.v(184)
    assign sha_core_block_read_data_next[34] = n305 ? xram_data_in[2] : sha_core_block[34];   // sha_top.v(184)
    assign sha_core_block_read_data_next[33] = n305 ? xram_data_in[1] : sha_core_block[33];   // sha_top.v(184)
    assign sha_core_block_read_data_next[32] = n305 ? xram_data_in[0] : sha_core_block[32];   // sha_top.v(184)
    nor (n318, n219, n218, n217, byte_counter[2], n215, byte_counter[0]) ;   // sha_top.v(185)
    assign sha_core_block_read_data_next[47] = n318 ? xram_data_in[7] : sha_core_block[47];   // sha_top.v(185)
    assign sha_core_block_read_data_next[46] = n318 ? xram_data_in[6] : sha_core_block[46];   // sha_top.v(185)
    assign sha_core_block_read_data_next[45] = n318 ? xram_data_in[5] : sha_core_block[45];   // sha_top.v(185)
    assign sha_core_block_read_data_next[44] = n318 ? xram_data_in[4] : sha_core_block[44];   // sha_top.v(185)
    assign sha_core_block_read_data_next[43] = n318 ? xram_data_in[3] : sha_core_block[43];   // sha_top.v(185)
    assign sha_core_block_read_data_next[42] = n318 ? xram_data_in[2] : sha_core_block[42];   // sha_top.v(185)
    assign sha_core_block_read_data_next[41] = n318 ? xram_data_in[1] : sha_core_block[41];   // sha_top.v(185)
    assign sha_core_block_read_data_next[40] = n318 ? xram_data_in[0] : sha_core_block[40];   // sha_top.v(185)
    nor (n331, n219, n218, n217, byte_counter[2], byte_counter[1], 
        n214) ;   // sha_top.v(186)
    assign sha_core_block_read_data_next[55] = n331 ? xram_data_in[7] : sha_core_block[55];   // sha_top.v(186)
    assign sha_core_block_read_data_next[54] = n331 ? xram_data_in[6] : sha_core_block[54];   // sha_top.v(186)
    assign sha_core_block_read_data_next[53] = n331 ? xram_data_in[5] : sha_core_block[53];   // sha_top.v(186)
    assign sha_core_block_read_data_next[52] = n331 ? xram_data_in[4] : sha_core_block[52];   // sha_top.v(186)
    assign sha_core_block_read_data_next[51] = n331 ? xram_data_in[3] : sha_core_block[51];   // sha_top.v(186)
    assign sha_core_block_read_data_next[50] = n331 ? xram_data_in[2] : sha_core_block[50];   // sha_top.v(186)
    assign sha_core_block_read_data_next[49] = n331 ? xram_data_in[1] : sha_core_block[49];   // sha_top.v(186)
    assign sha_core_block_read_data_next[48] = n331 ? xram_data_in[0] : sha_core_block[48];   // sha_top.v(186)
    nor (n343, n219, n218, n217, byte_counter[2], byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(187)
    assign sha_core_block_read_data_next[63] = n343 ? xram_data_in[7] : sha_core_block[63];   // sha_top.v(187)
    assign sha_core_block_read_data_next[62] = n343 ? xram_data_in[6] : sha_core_block[62];   // sha_top.v(187)
    assign sha_core_block_read_data_next[61] = n343 ? xram_data_in[5] : sha_core_block[61];   // sha_top.v(187)
    assign sha_core_block_read_data_next[60] = n343 ? xram_data_in[4] : sha_core_block[60];   // sha_top.v(187)
    assign sha_core_block_read_data_next[59] = n343 ? xram_data_in[3] : sha_core_block[59];   // sha_top.v(187)
    assign sha_core_block_read_data_next[58] = n343 ? xram_data_in[2] : sha_core_block[58];   // sha_top.v(187)
    assign sha_core_block_read_data_next[57] = n343 ? xram_data_in[1] : sha_core_block[57];   // sha_top.v(187)
    assign sha_core_block_read_data_next[56] = n343 ? xram_data_in[0] : sha_core_block[56];   // sha_top.v(187)
    nor (n357, n219, n218, byte_counter[3], n216, n215, n214) ;   // sha_top.v(188)
    assign sha_core_block_read_data_next[71] = n357 ? xram_data_in[7] : sha_core_block[71];   // sha_top.v(188)
    assign sha_core_block_read_data_next[70] = n357 ? xram_data_in[6] : sha_core_block[70];   // sha_top.v(188)
    assign sha_core_block_read_data_next[69] = n357 ? xram_data_in[5] : sha_core_block[69];   // sha_top.v(188)
    assign sha_core_block_read_data_next[68] = n357 ? xram_data_in[4] : sha_core_block[68];   // sha_top.v(188)
    assign sha_core_block_read_data_next[67] = n357 ? xram_data_in[3] : sha_core_block[67];   // sha_top.v(188)
    assign sha_core_block_read_data_next[66] = n357 ? xram_data_in[2] : sha_core_block[66];   // sha_top.v(188)
    assign sha_core_block_read_data_next[65] = n357 ? xram_data_in[1] : sha_core_block[65];   // sha_top.v(188)
    assign sha_core_block_read_data_next[64] = n357 ? xram_data_in[0] : sha_core_block[64];   // sha_top.v(188)
    nor (n370, n219, n218, byte_counter[3], n216, n215, byte_counter[0]) ;   // sha_top.v(189)
    assign sha_core_block_read_data_next[79] = n370 ? xram_data_in[7] : sha_core_block[79];   // sha_top.v(189)
    assign sha_core_block_read_data_next[78] = n370 ? xram_data_in[6] : sha_core_block[78];   // sha_top.v(189)
    assign sha_core_block_read_data_next[77] = n370 ? xram_data_in[5] : sha_core_block[77];   // sha_top.v(189)
    assign sha_core_block_read_data_next[76] = n370 ? xram_data_in[4] : sha_core_block[76];   // sha_top.v(189)
    assign sha_core_block_read_data_next[75] = n370 ? xram_data_in[3] : sha_core_block[75];   // sha_top.v(189)
    assign sha_core_block_read_data_next[74] = n370 ? xram_data_in[2] : sha_core_block[74];   // sha_top.v(189)
    assign sha_core_block_read_data_next[73] = n370 ? xram_data_in[1] : sha_core_block[73];   // sha_top.v(189)
    assign sha_core_block_read_data_next[72] = n370 ? xram_data_in[0] : sha_core_block[72];   // sha_top.v(189)
    nor (n383, n219, n218, byte_counter[3], n216, byte_counter[1], 
        n214) ;   // sha_top.v(190)
    assign sha_core_block_read_data_next[87] = n383 ? xram_data_in[7] : sha_core_block[87];   // sha_top.v(190)
    assign sha_core_block_read_data_next[86] = n383 ? xram_data_in[6] : sha_core_block[86];   // sha_top.v(190)
    assign sha_core_block_read_data_next[85] = n383 ? xram_data_in[5] : sha_core_block[85];   // sha_top.v(190)
    assign sha_core_block_read_data_next[84] = n383 ? xram_data_in[4] : sha_core_block[84];   // sha_top.v(190)
    assign sha_core_block_read_data_next[83] = n383 ? xram_data_in[3] : sha_core_block[83];   // sha_top.v(190)
    assign sha_core_block_read_data_next[82] = n383 ? xram_data_in[2] : sha_core_block[82];   // sha_top.v(190)
    assign sha_core_block_read_data_next[81] = n383 ? xram_data_in[1] : sha_core_block[81];   // sha_top.v(190)
    assign sha_core_block_read_data_next[80] = n383 ? xram_data_in[0] : sha_core_block[80];   // sha_top.v(190)
    nor (n395, n219, n218, byte_counter[3], n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(191)
    assign sha_core_block_read_data_next[95] = n395 ? xram_data_in[7] : sha_core_block[95];   // sha_top.v(191)
    assign sha_core_block_read_data_next[94] = n395 ? xram_data_in[6] : sha_core_block[94];   // sha_top.v(191)
    assign sha_core_block_read_data_next[93] = n395 ? xram_data_in[5] : sha_core_block[93];   // sha_top.v(191)
    assign sha_core_block_read_data_next[92] = n395 ? xram_data_in[4] : sha_core_block[92];   // sha_top.v(191)
    assign sha_core_block_read_data_next[91] = n395 ? xram_data_in[3] : sha_core_block[91];   // sha_top.v(191)
    assign sha_core_block_read_data_next[90] = n395 ? xram_data_in[2] : sha_core_block[90];   // sha_top.v(191)
    assign sha_core_block_read_data_next[89] = n395 ? xram_data_in[1] : sha_core_block[89];   // sha_top.v(191)
    assign sha_core_block_read_data_next[88] = n395 ? xram_data_in[0] : sha_core_block[88];   // sha_top.v(191)
    nor (n408, n219, n218, byte_counter[3], byte_counter[2], n215, 
        n214) ;   // sha_top.v(192)
    assign sha_core_block_read_data_next[103] = n408 ? xram_data_in[7] : sha_core_block[103];   // sha_top.v(192)
    assign sha_core_block_read_data_next[102] = n408 ? xram_data_in[6] : sha_core_block[102];   // sha_top.v(192)
    assign sha_core_block_read_data_next[101] = n408 ? xram_data_in[5] : sha_core_block[101];   // sha_top.v(192)
    assign sha_core_block_read_data_next[100] = n408 ? xram_data_in[4] : sha_core_block[100];   // sha_top.v(192)
    assign sha_core_block_read_data_next[99] = n408 ? xram_data_in[3] : sha_core_block[99];   // sha_top.v(192)
    assign sha_core_block_read_data_next[98] = n408 ? xram_data_in[2] : sha_core_block[98];   // sha_top.v(192)
    assign sha_core_block_read_data_next[97] = n408 ? xram_data_in[1] : sha_core_block[97];   // sha_top.v(192)
    assign sha_core_block_read_data_next[96] = n408 ? xram_data_in[0] : sha_core_block[96];   // sha_top.v(192)
    nor (n420, n219, n218, byte_counter[3], byte_counter[2], n215, 
        byte_counter[0]) ;   // sha_top.v(193)
    assign sha_core_block_read_data_next[111] = n420 ? xram_data_in[7] : sha_core_block[111];   // sha_top.v(193)
    assign sha_core_block_read_data_next[110] = n420 ? xram_data_in[6] : sha_core_block[110];   // sha_top.v(193)
    assign sha_core_block_read_data_next[109] = n420 ? xram_data_in[5] : sha_core_block[109];   // sha_top.v(193)
    assign sha_core_block_read_data_next[108] = n420 ? xram_data_in[4] : sha_core_block[108];   // sha_top.v(193)
    assign sha_core_block_read_data_next[107] = n420 ? xram_data_in[3] : sha_core_block[107];   // sha_top.v(193)
    assign sha_core_block_read_data_next[106] = n420 ? xram_data_in[2] : sha_core_block[106];   // sha_top.v(193)
    assign sha_core_block_read_data_next[105] = n420 ? xram_data_in[1] : sha_core_block[105];   // sha_top.v(193)
    assign sha_core_block_read_data_next[104] = n420 ? xram_data_in[0] : sha_core_block[104];   // sha_top.v(193)
    nor (n432, n219, n218, byte_counter[3], byte_counter[2], byte_counter[1], 
        n214) ;   // sha_top.v(194)
    assign sha_core_block_read_data_next[119] = n432 ? xram_data_in[7] : sha_core_block[119];   // sha_top.v(194)
    assign sha_core_block_read_data_next[118] = n432 ? xram_data_in[6] : sha_core_block[118];   // sha_top.v(194)
    assign sha_core_block_read_data_next[117] = n432 ? xram_data_in[5] : sha_core_block[117];   // sha_top.v(194)
    assign sha_core_block_read_data_next[116] = n432 ? xram_data_in[4] : sha_core_block[116];   // sha_top.v(194)
    assign sha_core_block_read_data_next[115] = n432 ? xram_data_in[3] : sha_core_block[115];   // sha_top.v(194)
    assign sha_core_block_read_data_next[114] = n432 ? xram_data_in[2] : sha_core_block[114];   // sha_top.v(194)
    assign sha_core_block_read_data_next[113] = n432 ? xram_data_in[1] : sha_core_block[113];   // sha_top.v(194)
    assign sha_core_block_read_data_next[112] = n432 ? xram_data_in[0] : sha_core_block[112];   // sha_top.v(194)
    nor (n443, n219, n218, byte_counter[3], byte_counter[2], byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(195)
    assign sha_core_block_read_data_next[127] = n443 ? xram_data_in[7] : sha_core_block[127];   // sha_top.v(195)
    assign sha_core_block_read_data_next[126] = n443 ? xram_data_in[6] : sha_core_block[126];   // sha_top.v(195)
    assign sha_core_block_read_data_next[125] = n443 ? xram_data_in[5] : sha_core_block[125];   // sha_top.v(195)
    assign sha_core_block_read_data_next[124] = n443 ? xram_data_in[4] : sha_core_block[124];   // sha_top.v(195)
    assign sha_core_block_read_data_next[123] = n443 ? xram_data_in[3] : sha_core_block[123];   // sha_top.v(195)
    assign sha_core_block_read_data_next[122] = n443 ? xram_data_in[2] : sha_core_block[122];   // sha_top.v(195)
    assign sha_core_block_read_data_next[121] = n443 ? xram_data_in[1] : sha_core_block[121];   // sha_top.v(195)
    assign sha_core_block_read_data_next[120] = n443 ? xram_data_in[0] : sha_core_block[120];   // sha_top.v(195)
    nor (n457, n219, byte_counter[4], n217, n216, n215, n214) ;   // sha_top.v(196)
    assign sha_core_block_read_data_next[135] = n457 ? xram_data_in[7] : sha_core_block[135];   // sha_top.v(196)
    assign sha_core_block_read_data_next[134] = n457 ? xram_data_in[6] : sha_core_block[134];   // sha_top.v(196)
    assign sha_core_block_read_data_next[133] = n457 ? xram_data_in[5] : sha_core_block[133];   // sha_top.v(196)
    assign sha_core_block_read_data_next[132] = n457 ? xram_data_in[4] : sha_core_block[132];   // sha_top.v(196)
    assign sha_core_block_read_data_next[131] = n457 ? xram_data_in[3] : sha_core_block[131];   // sha_top.v(196)
    assign sha_core_block_read_data_next[130] = n457 ? xram_data_in[2] : sha_core_block[130];   // sha_top.v(196)
    assign sha_core_block_read_data_next[129] = n457 ? xram_data_in[1] : sha_core_block[129];   // sha_top.v(196)
    assign sha_core_block_read_data_next[128] = n457 ? xram_data_in[0] : sha_core_block[128];   // sha_top.v(196)
    nor (n470, n219, byte_counter[4], n217, n216, n215, byte_counter[0]) ;   // sha_top.v(197)
    assign sha_core_block_read_data_next[143] = n470 ? xram_data_in[7] : sha_core_block[143];   // sha_top.v(197)
    assign sha_core_block_read_data_next[142] = n470 ? xram_data_in[6] : sha_core_block[142];   // sha_top.v(197)
    assign sha_core_block_read_data_next[141] = n470 ? xram_data_in[5] : sha_core_block[141];   // sha_top.v(197)
    assign sha_core_block_read_data_next[140] = n470 ? xram_data_in[4] : sha_core_block[140];   // sha_top.v(197)
    assign sha_core_block_read_data_next[139] = n470 ? xram_data_in[3] : sha_core_block[139];   // sha_top.v(197)
    assign sha_core_block_read_data_next[138] = n470 ? xram_data_in[2] : sha_core_block[138];   // sha_top.v(197)
    assign sha_core_block_read_data_next[137] = n470 ? xram_data_in[1] : sha_core_block[137];   // sha_top.v(197)
    assign sha_core_block_read_data_next[136] = n470 ? xram_data_in[0] : sha_core_block[136];   // sha_top.v(197)
    nor (n483, n219, byte_counter[4], n217, n216, byte_counter[1], 
        n214) ;   // sha_top.v(198)
    assign sha_core_block_read_data_next[151] = n483 ? xram_data_in[7] : sha_core_block[151];   // sha_top.v(198)
    assign sha_core_block_read_data_next[150] = n483 ? xram_data_in[6] : sha_core_block[150];   // sha_top.v(198)
    assign sha_core_block_read_data_next[149] = n483 ? xram_data_in[5] : sha_core_block[149];   // sha_top.v(198)
    assign sha_core_block_read_data_next[148] = n483 ? xram_data_in[4] : sha_core_block[148];   // sha_top.v(198)
    assign sha_core_block_read_data_next[147] = n483 ? xram_data_in[3] : sha_core_block[147];   // sha_top.v(198)
    assign sha_core_block_read_data_next[146] = n483 ? xram_data_in[2] : sha_core_block[146];   // sha_top.v(198)
    assign sha_core_block_read_data_next[145] = n483 ? xram_data_in[1] : sha_core_block[145];   // sha_top.v(198)
    assign sha_core_block_read_data_next[144] = n483 ? xram_data_in[0] : sha_core_block[144];   // sha_top.v(198)
    nor (n495, n219, byte_counter[4], n217, n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(199)
    assign sha_core_block_read_data_next[159] = n495 ? xram_data_in[7] : sha_core_block[159];   // sha_top.v(199)
    assign sha_core_block_read_data_next[158] = n495 ? xram_data_in[6] : sha_core_block[158];   // sha_top.v(199)
    assign sha_core_block_read_data_next[157] = n495 ? xram_data_in[5] : sha_core_block[157];   // sha_top.v(199)
    assign sha_core_block_read_data_next[156] = n495 ? xram_data_in[4] : sha_core_block[156];   // sha_top.v(199)
    assign sha_core_block_read_data_next[155] = n495 ? xram_data_in[3] : sha_core_block[155];   // sha_top.v(199)
    assign sha_core_block_read_data_next[154] = n495 ? xram_data_in[2] : sha_core_block[154];   // sha_top.v(199)
    assign sha_core_block_read_data_next[153] = n495 ? xram_data_in[1] : sha_core_block[153];   // sha_top.v(199)
    assign sha_core_block_read_data_next[152] = n495 ? xram_data_in[0] : sha_core_block[152];   // sha_top.v(199)
    nor (n508, n219, byte_counter[4], n217, byte_counter[2], n215, 
        n214) ;   // sha_top.v(200)
    assign sha_core_block_read_data_next[167] = n508 ? xram_data_in[7] : sha_core_block[167];   // sha_top.v(200)
    assign sha_core_block_read_data_next[166] = n508 ? xram_data_in[6] : sha_core_block[166];   // sha_top.v(200)
    assign sha_core_block_read_data_next[165] = n508 ? xram_data_in[5] : sha_core_block[165];   // sha_top.v(200)
    assign sha_core_block_read_data_next[164] = n508 ? xram_data_in[4] : sha_core_block[164];   // sha_top.v(200)
    assign sha_core_block_read_data_next[163] = n508 ? xram_data_in[3] : sha_core_block[163];   // sha_top.v(200)
    assign sha_core_block_read_data_next[162] = n508 ? xram_data_in[2] : sha_core_block[162];   // sha_top.v(200)
    assign sha_core_block_read_data_next[161] = n508 ? xram_data_in[1] : sha_core_block[161];   // sha_top.v(200)
    assign sha_core_block_read_data_next[160] = n508 ? xram_data_in[0] : sha_core_block[160];   // sha_top.v(200)
    nor (n520, n219, byte_counter[4], n217, byte_counter[2], n215, 
        byte_counter[0]) ;   // sha_top.v(201)
    assign sha_core_block_read_data_next[175] = n520 ? xram_data_in[7] : sha_core_block[175];   // sha_top.v(201)
    assign sha_core_block_read_data_next[174] = n520 ? xram_data_in[6] : sha_core_block[174];   // sha_top.v(201)
    assign sha_core_block_read_data_next[173] = n520 ? xram_data_in[5] : sha_core_block[173];   // sha_top.v(201)
    assign sha_core_block_read_data_next[172] = n520 ? xram_data_in[4] : sha_core_block[172];   // sha_top.v(201)
    assign sha_core_block_read_data_next[171] = n520 ? xram_data_in[3] : sha_core_block[171];   // sha_top.v(201)
    assign sha_core_block_read_data_next[170] = n520 ? xram_data_in[2] : sha_core_block[170];   // sha_top.v(201)
    assign sha_core_block_read_data_next[169] = n520 ? xram_data_in[1] : sha_core_block[169];   // sha_top.v(201)
    assign sha_core_block_read_data_next[168] = n520 ? xram_data_in[0] : sha_core_block[168];   // sha_top.v(201)
    nor (n532, n219, byte_counter[4], n217, byte_counter[2], byte_counter[1], 
        n214) ;   // sha_top.v(202)
    assign sha_core_block_read_data_next[183] = n532 ? xram_data_in[7] : sha_core_block[183];   // sha_top.v(202)
    assign sha_core_block_read_data_next[182] = n532 ? xram_data_in[6] : sha_core_block[182];   // sha_top.v(202)
    assign sha_core_block_read_data_next[181] = n532 ? xram_data_in[5] : sha_core_block[181];   // sha_top.v(202)
    assign sha_core_block_read_data_next[180] = n532 ? xram_data_in[4] : sha_core_block[180];   // sha_top.v(202)
    assign sha_core_block_read_data_next[179] = n532 ? xram_data_in[3] : sha_core_block[179];   // sha_top.v(202)
    assign sha_core_block_read_data_next[178] = n532 ? xram_data_in[2] : sha_core_block[178];   // sha_top.v(202)
    assign sha_core_block_read_data_next[177] = n532 ? xram_data_in[1] : sha_core_block[177];   // sha_top.v(202)
    assign sha_core_block_read_data_next[176] = n532 ? xram_data_in[0] : sha_core_block[176];   // sha_top.v(202)
    nor (n543, n219, byte_counter[4], n217, byte_counter[2], byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(203)
    assign sha_core_block_read_data_next[191] = n543 ? xram_data_in[7] : sha_core_block[191];   // sha_top.v(203)
    assign sha_core_block_read_data_next[190] = n543 ? xram_data_in[6] : sha_core_block[190];   // sha_top.v(203)
    assign sha_core_block_read_data_next[189] = n543 ? xram_data_in[5] : sha_core_block[189];   // sha_top.v(203)
    assign sha_core_block_read_data_next[188] = n543 ? xram_data_in[4] : sha_core_block[188];   // sha_top.v(203)
    assign sha_core_block_read_data_next[187] = n543 ? xram_data_in[3] : sha_core_block[187];   // sha_top.v(203)
    assign sha_core_block_read_data_next[186] = n543 ? xram_data_in[2] : sha_core_block[186];   // sha_top.v(203)
    assign sha_core_block_read_data_next[185] = n543 ? xram_data_in[1] : sha_core_block[185];   // sha_top.v(203)
    assign sha_core_block_read_data_next[184] = n543 ? xram_data_in[0] : sha_core_block[184];   // sha_top.v(203)
    nor (n556, n219, byte_counter[4], byte_counter[3], n216, n215, 
        n214) ;   // sha_top.v(204)
    assign sha_core_block_read_data_next[199] = n556 ? xram_data_in[7] : sha_core_block[199];   // sha_top.v(204)
    assign sha_core_block_read_data_next[198] = n556 ? xram_data_in[6] : sha_core_block[198];   // sha_top.v(204)
    assign sha_core_block_read_data_next[197] = n556 ? xram_data_in[5] : sha_core_block[197];   // sha_top.v(204)
    assign sha_core_block_read_data_next[196] = n556 ? xram_data_in[4] : sha_core_block[196];   // sha_top.v(204)
    assign sha_core_block_read_data_next[195] = n556 ? xram_data_in[3] : sha_core_block[195];   // sha_top.v(204)
    assign sha_core_block_read_data_next[194] = n556 ? xram_data_in[2] : sha_core_block[194];   // sha_top.v(204)
    assign sha_core_block_read_data_next[193] = n556 ? xram_data_in[1] : sha_core_block[193];   // sha_top.v(204)
    assign sha_core_block_read_data_next[192] = n556 ? xram_data_in[0] : sha_core_block[192];   // sha_top.v(204)
    nor (n568, n219, byte_counter[4], byte_counter[3], n216, n215, 
        byte_counter[0]) ;   // sha_top.v(205)
    assign sha_core_block_read_data_next[207] = n568 ? xram_data_in[7] : sha_core_block[207];   // sha_top.v(205)
    assign sha_core_block_read_data_next[206] = n568 ? xram_data_in[6] : sha_core_block[206];   // sha_top.v(205)
    assign sha_core_block_read_data_next[205] = n568 ? xram_data_in[5] : sha_core_block[205];   // sha_top.v(205)
    assign sha_core_block_read_data_next[204] = n568 ? xram_data_in[4] : sha_core_block[204];   // sha_top.v(205)
    assign sha_core_block_read_data_next[203] = n568 ? xram_data_in[3] : sha_core_block[203];   // sha_top.v(205)
    assign sha_core_block_read_data_next[202] = n568 ? xram_data_in[2] : sha_core_block[202];   // sha_top.v(205)
    assign sha_core_block_read_data_next[201] = n568 ? xram_data_in[1] : sha_core_block[201];   // sha_top.v(205)
    assign sha_core_block_read_data_next[200] = n568 ? xram_data_in[0] : sha_core_block[200];   // sha_top.v(205)
    nor (n580, n219, byte_counter[4], byte_counter[3], n216, byte_counter[1], 
        n214) ;   // sha_top.v(206)
    assign sha_core_block_read_data_next[215] = n580 ? xram_data_in[7] : sha_core_block[215];   // sha_top.v(206)
    assign sha_core_block_read_data_next[214] = n580 ? xram_data_in[6] : sha_core_block[214];   // sha_top.v(206)
    assign sha_core_block_read_data_next[213] = n580 ? xram_data_in[5] : sha_core_block[213];   // sha_top.v(206)
    assign sha_core_block_read_data_next[212] = n580 ? xram_data_in[4] : sha_core_block[212];   // sha_top.v(206)
    assign sha_core_block_read_data_next[211] = n580 ? xram_data_in[3] : sha_core_block[211];   // sha_top.v(206)
    assign sha_core_block_read_data_next[210] = n580 ? xram_data_in[2] : sha_core_block[210];   // sha_top.v(206)
    assign sha_core_block_read_data_next[209] = n580 ? xram_data_in[1] : sha_core_block[209];   // sha_top.v(206)
    assign sha_core_block_read_data_next[208] = n580 ? xram_data_in[0] : sha_core_block[208];   // sha_top.v(206)
    nor (n591, n219, byte_counter[4], byte_counter[3], n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(207)
    assign sha_core_block_read_data_next[223] = n591 ? xram_data_in[7] : sha_core_block[223];   // sha_top.v(207)
    assign sha_core_block_read_data_next[222] = n591 ? xram_data_in[6] : sha_core_block[222];   // sha_top.v(207)
    assign sha_core_block_read_data_next[221] = n591 ? xram_data_in[5] : sha_core_block[221];   // sha_top.v(207)
    assign sha_core_block_read_data_next[220] = n591 ? xram_data_in[4] : sha_core_block[220];   // sha_top.v(207)
    assign sha_core_block_read_data_next[219] = n591 ? xram_data_in[3] : sha_core_block[219];   // sha_top.v(207)
    assign sha_core_block_read_data_next[218] = n591 ? xram_data_in[2] : sha_core_block[218];   // sha_top.v(207)
    assign sha_core_block_read_data_next[217] = n591 ? xram_data_in[1] : sha_core_block[217];   // sha_top.v(207)
    assign sha_core_block_read_data_next[216] = n591 ? xram_data_in[0] : sha_core_block[216];   // sha_top.v(207)
    nor (n603, n219, byte_counter[4], byte_counter[3], byte_counter[2], 
        n215, n214) ;   // sha_top.v(208)
    assign sha_core_block_read_data_next[231] = n603 ? xram_data_in[7] : sha_core_block[231];   // sha_top.v(208)
    assign sha_core_block_read_data_next[230] = n603 ? xram_data_in[6] : sha_core_block[230];   // sha_top.v(208)
    assign sha_core_block_read_data_next[229] = n603 ? xram_data_in[5] : sha_core_block[229];   // sha_top.v(208)
    assign sha_core_block_read_data_next[228] = n603 ? xram_data_in[4] : sha_core_block[228];   // sha_top.v(208)
    assign sha_core_block_read_data_next[227] = n603 ? xram_data_in[3] : sha_core_block[227];   // sha_top.v(208)
    assign sha_core_block_read_data_next[226] = n603 ? xram_data_in[2] : sha_core_block[226];   // sha_top.v(208)
    assign sha_core_block_read_data_next[225] = n603 ? xram_data_in[1] : sha_core_block[225];   // sha_top.v(208)
    assign sha_core_block_read_data_next[224] = n603 ? xram_data_in[0] : sha_core_block[224];   // sha_top.v(208)
    nor (n614, n219, byte_counter[4], byte_counter[3], byte_counter[2], 
        n215, byte_counter[0]) ;   // sha_top.v(209)
    assign sha_core_block_read_data_next[239] = n614 ? xram_data_in[7] : sha_core_block[239];   // sha_top.v(209)
    assign sha_core_block_read_data_next[238] = n614 ? xram_data_in[6] : sha_core_block[238];   // sha_top.v(209)
    assign sha_core_block_read_data_next[237] = n614 ? xram_data_in[5] : sha_core_block[237];   // sha_top.v(209)
    assign sha_core_block_read_data_next[236] = n614 ? xram_data_in[4] : sha_core_block[236];   // sha_top.v(209)
    assign sha_core_block_read_data_next[235] = n614 ? xram_data_in[3] : sha_core_block[235];   // sha_top.v(209)
    assign sha_core_block_read_data_next[234] = n614 ? xram_data_in[2] : sha_core_block[234];   // sha_top.v(209)
    assign sha_core_block_read_data_next[233] = n614 ? xram_data_in[1] : sha_core_block[233];   // sha_top.v(209)
    assign sha_core_block_read_data_next[232] = n614 ? xram_data_in[0] : sha_core_block[232];   // sha_top.v(209)
    nor (n625, n219, byte_counter[4], byte_counter[3], byte_counter[2], 
        byte_counter[1], n214) ;   // sha_top.v(210)
    assign sha_core_block_read_data_next[247] = n625 ? xram_data_in[7] : sha_core_block[247];   // sha_top.v(210)
    assign sha_core_block_read_data_next[246] = n625 ? xram_data_in[6] : sha_core_block[246];   // sha_top.v(210)
    assign sha_core_block_read_data_next[245] = n625 ? xram_data_in[5] : sha_core_block[245];   // sha_top.v(210)
    assign sha_core_block_read_data_next[244] = n625 ? xram_data_in[4] : sha_core_block[244];   // sha_top.v(210)
    assign sha_core_block_read_data_next[243] = n625 ? xram_data_in[3] : sha_core_block[243];   // sha_top.v(210)
    assign sha_core_block_read_data_next[242] = n625 ? xram_data_in[2] : sha_core_block[242];   // sha_top.v(210)
    assign sha_core_block_read_data_next[241] = n625 ? xram_data_in[1] : sha_core_block[241];   // sha_top.v(210)
    assign sha_core_block_read_data_next[240] = n625 ? xram_data_in[0] : sha_core_block[240];   // sha_top.v(210)
    nor (n635, n219, byte_counter[4], byte_counter[3], byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // sha_top.v(211)
    assign sha_core_block_read_data_next[255] = n635 ? xram_data_in[7] : sha_core_block[255];   // sha_top.v(211)
    assign sha_core_block_read_data_next[254] = n635 ? xram_data_in[6] : sha_core_block[254];   // sha_top.v(211)
    assign sha_core_block_read_data_next[253] = n635 ? xram_data_in[5] : sha_core_block[253];   // sha_top.v(211)
    assign sha_core_block_read_data_next[252] = n635 ? xram_data_in[4] : sha_core_block[252];   // sha_top.v(211)
    assign sha_core_block_read_data_next[251] = n635 ? xram_data_in[3] : sha_core_block[251];   // sha_top.v(211)
    assign sha_core_block_read_data_next[250] = n635 ? xram_data_in[2] : sha_core_block[250];   // sha_top.v(211)
    assign sha_core_block_read_data_next[249] = n635 ? xram_data_in[1] : sha_core_block[249];   // sha_top.v(211)
    assign sha_core_block_read_data_next[248] = n635 ? xram_data_in[0] : sha_core_block[248];   // sha_top.v(211)
    nor (n649, byte_counter[5], n218, n217, n216, n215, n214) ;   // sha_top.v(212)
    assign sha_core_block_read_data_next[263] = n649 ? xram_data_in[7] : sha_core_block[263];   // sha_top.v(212)
    assign sha_core_block_read_data_next[262] = n649 ? xram_data_in[6] : sha_core_block[262];   // sha_top.v(212)
    assign sha_core_block_read_data_next[261] = n649 ? xram_data_in[5] : sha_core_block[261];   // sha_top.v(212)
    assign sha_core_block_read_data_next[260] = n649 ? xram_data_in[4] : sha_core_block[260];   // sha_top.v(212)
    assign sha_core_block_read_data_next[259] = n649 ? xram_data_in[3] : sha_core_block[259];   // sha_top.v(212)
    assign sha_core_block_read_data_next[258] = n649 ? xram_data_in[2] : sha_core_block[258];   // sha_top.v(212)
    assign sha_core_block_read_data_next[257] = n649 ? xram_data_in[1] : sha_core_block[257];   // sha_top.v(212)
    assign sha_core_block_read_data_next[256] = n649 ? xram_data_in[0] : sha_core_block[256];   // sha_top.v(212)
    nor (n662, byte_counter[5], n218, n217, n216, n215, byte_counter[0]) ;   // sha_top.v(213)
    assign sha_core_block_read_data_next[271] = n662 ? xram_data_in[7] : sha_core_block[271];   // sha_top.v(213)
    assign sha_core_block_read_data_next[270] = n662 ? xram_data_in[6] : sha_core_block[270];   // sha_top.v(213)
    assign sha_core_block_read_data_next[269] = n662 ? xram_data_in[5] : sha_core_block[269];   // sha_top.v(213)
    assign sha_core_block_read_data_next[268] = n662 ? xram_data_in[4] : sha_core_block[268];   // sha_top.v(213)
    assign sha_core_block_read_data_next[267] = n662 ? xram_data_in[3] : sha_core_block[267];   // sha_top.v(213)
    assign sha_core_block_read_data_next[266] = n662 ? xram_data_in[2] : sha_core_block[266];   // sha_top.v(213)
    assign sha_core_block_read_data_next[265] = n662 ? xram_data_in[1] : sha_core_block[265];   // sha_top.v(213)
    assign sha_core_block_read_data_next[264] = n662 ? xram_data_in[0] : sha_core_block[264];   // sha_top.v(213)
    nor (n675, byte_counter[5], n218, n217, n216, byte_counter[1], 
        n214) ;   // sha_top.v(214)
    assign sha_core_block_read_data_next[279] = n675 ? xram_data_in[7] : sha_core_block[279];   // sha_top.v(214)
    assign sha_core_block_read_data_next[278] = n675 ? xram_data_in[6] : sha_core_block[278];   // sha_top.v(214)
    assign sha_core_block_read_data_next[277] = n675 ? xram_data_in[5] : sha_core_block[277];   // sha_top.v(214)
    assign sha_core_block_read_data_next[276] = n675 ? xram_data_in[4] : sha_core_block[276];   // sha_top.v(214)
    assign sha_core_block_read_data_next[275] = n675 ? xram_data_in[3] : sha_core_block[275];   // sha_top.v(214)
    assign sha_core_block_read_data_next[274] = n675 ? xram_data_in[2] : sha_core_block[274];   // sha_top.v(214)
    assign sha_core_block_read_data_next[273] = n675 ? xram_data_in[1] : sha_core_block[273];   // sha_top.v(214)
    assign sha_core_block_read_data_next[272] = n675 ? xram_data_in[0] : sha_core_block[272];   // sha_top.v(214)
    nor (n687, byte_counter[5], n218, n217, n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(215)
    assign sha_core_block_read_data_next[287] = n687 ? xram_data_in[7] : sha_core_block[287];   // sha_top.v(215)
    assign sha_core_block_read_data_next[286] = n687 ? xram_data_in[6] : sha_core_block[286];   // sha_top.v(215)
    assign sha_core_block_read_data_next[285] = n687 ? xram_data_in[5] : sha_core_block[285];   // sha_top.v(215)
    assign sha_core_block_read_data_next[284] = n687 ? xram_data_in[4] : sha_core_block[284];   // sha_top.v(215)
    assign sha_core_block_read_data_next[283] = n687 ? xram_data_in[3] : sha_core_block[283];   // sha_top.v(215)
    assign sha_core_block_read_data_next[282] = n687 ? xram_data_in[2] : sha_core_block[282];   // sha_top.v(215)
    assign sha_core_block_read_data_next[281] = n687 ? xram_data_in[1] : sha_core_block[281];   // sha_top.v(215)
    assign sha_core_block_read_data_next[280] = n687 ? xram_data_in[0] : sha_core_block[280];   // sha_top.v(215)
    nor (n700, byte_counter[5], n218, n217, byte_counter[2], n215, 
        n214) ;   // sha_top.v(216)
    assign sha_core_block_read_data_next[295] = n700 ? xram_data_in[7] : sha_core_block[295];   // sha_top.v(216)
    assign sha_core_block_read_data_next[294] = n700 ? xram_data_in[6] : sha_core_block[294];   // sha_top.v(216)
    assign sha_core_block_read_data_next[293] = n700 ? xram_data_in[5] : sha_core_block[293];   // sha_top.v(216)
    assign sha_core_block_read_data_next[292] = n700 ? xram_data_in[4] : sha_core_block[292];   // sha_top.v(216)
    assign sha_core_block_read_data_next[291] = n700 ? xram_data_in[3] : sha_core_block[291];   // sha_top.v(216)
    assign sha_core_block_read_data_next[290] = n700 ? xram_data_in[2] : sha_core_block[290];   // sha_top.v(216)
    assign sha_core_block_read_data_next[289] = n700 ? xram_data_in[1] : sha_core_block[289];   // sha_top.v(216)
    assign sha_core_block_read_data_next[288] = n700 ? xram_data_in[0] : sha_core_block[288];   // sha_top.v(216)
    nor (n712, byte_counter[5], n218, n217, byte_counter[2], n215, 
        byte_counter[0]) ;   // sha_top.v(217)
    assign sha_core_block_read_data_next[303] = n712 ? xram_data_in[7] : sha_core_block[303];   // sha_top.v(217)
    assign sha_core_block_read_data_next[302] = n712 ? xram_data_in[6] : sha_core_block[302];   // sha_top.v(217)
    assign sha_core_block_read_data_next[301] = n712 ? xram_data_in[5] : sha_core_block[301];   // sha_top.v(217)
    assign sha_core_block_read_data_next[300] = n712 ? xram_data_in[4] : sha_core_block[300];   // sha_top.v(217)
    assign sha_core_block_read_data_next[299] = n712 ? xram_data_in[3] : sha_core_block[299];   // sha_top.v(217)
    assign sha_core_block_read_data_next[298] = n712 ? xram_data_in[2] : sha_core_block[298];   // sha_top.v(217)
    assign sha_core_block_read_data_next[297] = n712 ? xram_data_in[1] : sha_core_block[297];   // sha_top.v(217)
    assign sha_core_block_read_data_next[296] = n712 ? xram_data_in[0] : sha_core_block[296];   // sha_top.v(217)
    nor (n724, byte_counter[5], n218, n217, byte_counter[2], byte_counter[1], 
        n214) ;   // sha_top.v(218)
    assign sha_core_block_read_data_next[311] = n724 ? xram_data_in[7] : sha_core_block[311];   // sha_top.v(218)
    assign sha_core_block_read_data_next[310] = n724 ? xram_data_in[6] : sha_core_block[310];   // sha_top.v(218)
    assign sha_core_block_read_data_next[309] = n724 ? xram_data_in[5] : sha_core_block[309];   // sha_top.v(218)
    assign sha_core_block_read_data_next[308] = n724 ? xram_data_in[4] : sha_core_block[308];   // sha_top.v(218)
    assign sha_core_block_read_data_next[307] = n724 ? xram_data_in[3] : sha_core_block[307];   // sha_top.v(218)
    assign sha_core_block_read_data_next[306] = n724 ? xram_data_in[2] : sha_core_block[306];   // sha_top.v(218)
    assign sha_core_block_read_data_next[305] = n724 ? xram_data_in[1] : sha_core_block[305];   // sha_top.v(218)
    assign sha_core_block_read_data_next[304] = n724 ? xram_data_in[0] : sha_core_block[304];   // sha_top.v(218)
    nor (n735, byte_counter[5], n218, n217, byte_counter[2], byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(219)
    assign sha_core_block_read_data_next[319] = n735 ? xram_data_in[7] : sha_core_block[319];   // sha_top.v(219)
    assign sha_core_block_read_data_next[318] = n735 ? xram_data_in[6] : sha_core_block[318];   // sha_top.v(219)
    assign sha_core_block_read_data_next[317] = n735 ? xram_data_in[5] : sha_core_block[317];   // sha_top.v(219)
    assign sha_core_block_read_data_next[316] = n735 ? xram_data_in[4] : sha_core_block[316];   // sha_top.v(219)
    assign sha_core_block_read_data_next[315] = n735 ? xram_data_in[3] : sha_core_block[315];   // sha_top.v(219)
    assign sha_core_block_read_data_next[314] = n735 ? xram_data_in[2] : sha_core_block[314];   // sha_top.v(219)
    assign sha_core_block_read_data_next[313] = n735 ? xram_data_in[1] : sha_core_block[313];   // sha_top.v(219)
    assign sha_core_block_read_data_next[312] = n735 ? xram_data_in[0] : sha_core_block[312];   // sha_top.v(219)
    nor (n748, byte_counter[5], n218, byte_counter[3], n216, n215, 
        n214) ;   // sha_top.v(220)
    assign sha_core_block_read_data_next[327] = n748 ? xram_data_in[7] : sha_core_block[327];   // sha_top.v(220)
    assign sha_core_block_read_data_next[326] = n748 ? xram_data_in[6] : sha_core_block[326];   // sha_top.v(220)
    assign sha_core_block_read_data_next[325] = n748 ? xram_data_in[5] : sha_core_block[325];   // sha_top.v(220)
    assign sha_core_block_read_data_next[324] = n748 ? xram_data_in[4] : sha_core_block[324];   // sha_top.v(220)
    assign sha_core_block_read_data_next[323] = n748 ? xram_data_in[3] : sha_core_block[323];   // sha_top.v(220)
    assign sha_core_block_read_data_next[322] = n748 ? xram_data_in[2] : sha_core_block[322];   // sha_top.v(220)
    assign sha_core_block_read_data_next[321] = n748 ? xram_data_in[1] : sha_core_block[321];   // sha_top.v(220)
    assign sha_core_block_read_data_next[320] = n748 ? xram_data_in[0] : sha_core_block[320];   // sha_top.v(220)
    nor (n760, byte_counter[5], n218, byte_counter[3], n216, n215, 
        byte_counter[0]) ;   // sha_top.v(221)
    assign sha_core_block_read_data_next[335] = n760 ? xram_data_in[7] : sha_core_block[335];   // sha_top.v(221)
    assign sha_core_block_read_data_next[334] = n760 ? xram_data_in[6] : sha_core_block[334];   // sha_top.v(221)
    assign sha_core_block_read_data_next[333] = n760 ? xram_data_in[5] : sha_core_block[333];   // sha_top.v(221)
    assign sha_core_block_read_data_next[332] = n760 ? xram_data_in[4] : sha_core_block[332];   // sha_top.v(221)
    assign sha_core_block_read_data_next[331] = n760 ? xram_data_in[3] : sha_core_block[331];   // sha_top.v(221)
    assign sha_core_block_read_data_next[330] = n760 ? xram_data_in[2] : sha_core_block[330];   // sha_top.v(221)
    assign sha_core_block_read_data_next[329] = n760 ? xram_data_in[1] : sha_core_block[329];   // sha_top.v(221)
    assign sha_core_block_read_data_next[328] = n760 ? xram_data_in[0] : sha_core_block[328];   // sha_top.v(221)
    nor (n772, byte_counter[5], n218, byte_counter[3], n216, byte_counter[1], 
        n214) ;   // sha_top.v(222)
    assign sha_core_block_read_data_next[343] = n772 ? xram_data_in[7] : sha_core_block[343];   // sha_top.v(222)
    assign sha_core_block_read_data_next[342] = n772 ? xram_data_in[6] : sha_core_block[342];   // sha_top.v(222)
    assign sha_core_block_read_data_next[341] = n772 ? xram_data_in[5] : sha_core_block[341];   // sha_top.v(222)
    assign sha_core_block_read_data_next[340] = n772 ? xram_data_in[4] : sha_core_block[340];   // sha_top.v(222)
    assign sha_core_block_read_data_next[339] = n772 ? xram_data_in[3] : sha_core_block[339];   // sha_top.v(222)
    assign sha_core_block_read_data_next[338] = n772 ? xram_data_in[2] : sha_core_block[338];   // sha_top.v(222)
    assign sha_core_block_read_data_next[337] = n772 ? xram_data_in[1] : sha_core_block[337];   // sha_top.v(222)
    assign sha_core_block_read_data_next[336] = n772 ? xram_data_in[0] : sha_core_block[336];   // sha_top.v(222)
    nor (n783, byte_counter[5], n218, byte_counter[3], n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(223)
    assign sha_core_block_read_data_next[351] = n783 ? xram_data_in[7] : sha_core_block[351];   // sha_top.v(223)
    assign sha_core_block_read_data_next[350] = n783 ? xram_data_in[6] : sha_core_block[350];   // sha_top.v(223)
    assign sha_core_block_read_data_next[349] = n783 ? xram_data_in[5] : sha_core_block[349];   // sha_top.v(223)
    assign sha_core_block_read_data_next[348] = n783 ? xram_data_in[4] : sha_core_block[348];   // sha_top.v(223)
    assign sha_core_block_read_data_next[347] = n783 ? xram_data_in[3] : sha_core_block[347];   // sha_top.v(223)
    assign sha_core_block_read_data_next[346] = n783 ? xram_data_in[2] : sha_core_block[346];   // sha_top.v(223)
    assign sha_core_block_read_data_next[345] = n783 ? xram_data_in[1] : sha_core_block[345];   // sha_top.v(223)
    assign sha_core_block_read_data_next[344] = n783 ? xram_data_in[0] : sha_core_block[344];   // sha_top.v(223)
    nor (writing_last_byte, byte_counter[5], n218, byte_counter[3], 
        byte_counter[2], n215, n214) ;   // sha_top.v(224)
    assign sha_core_block_read_data_next[359] = writing_last_byte ? xram_data_in[7] : sha_core_block[359];   // sha_top.v(224)
    assign sha_core_block_read_data_next[358] = writing_last_byte ? xram_data_in[6] : sha_core_block[358];   // sha_top.v(224)
    assign sha_core_block_read_data_next[357] = writing_last_byte ? xram_data_in[5] : sha_core_block[357];   // sha_top.v(224)
    assign sha_core_block_read_data_next[356] = writing_last_byte ? xram_data_in[4] : sha_core_block[356];   // sha_top.v(224)
    assign sha_core_block_read_data_next[355] = writing_last_byte ? xram_data_in[3] : sha_core_block[355];   // sha_top.v(224)
    assign sha_core_block_read_data_next[354] = writing_last_byte ? xram_data_in[2] : sha_core_block[354];   // sha_top.v(224)
    assign sha_core_block_read_data_next[353] = writing_last_byte ? xram_data_in[1] : sha_core_block[353];   // sha_top.v(224)
    assign sha_core_block_read_data_next[352] = writing_last_byte ? xram_data_in[0] : sha_core_block[352];   // sha_top.v(224)
    nor (n806, byte_counter[5], n218, byte_counter[3], byte_counter[2], 
        n215, byte_counter[0]) ;   // sha_top.v(225)
    assign sha_core_block_read_data_next[367] = n806 ? xram_data_in[7] : sha_core_block[367];   // sha_top.v(225)
    assign sha_core_block_read_data_next[366] = n806 ? xram_data_in[6] : sha_core_block[366];   // sha_top.v(225)
    assign sha_core_block_read_data_next[365] = n806 ? xram_data_in[5] : sha_core_block[365];   // sha_top.v(225)
    assign sha_core_block_read_data_next[364] = n806 ? xram_data_in[4] : sha_core_block[364];   // sha_top.v(225)
    assign sha_core_block_read_data_next[363] = n806 ? xram_data_in[3] : sha_core_block[363];   // sha_top.v(225)
    assign sha_core_block_read_data_next[362] = n806 ? xram_data_in[2] : sha_core_block[362];   // sha_top.v(225)
    assign sha_core_block_read_data_next[361] = n806 ? xram_data_in[1] : sha_core_block[361];   // sha_top.v(225)
    assign sha_core_block_read_data_next[360] = n806 ? xram_data_in[0] : sha_core_block[360];   // sha_top.v(225)
    nor (n817, byte_counter[5], n218, byte_counter[3], byte_counter[2], 
        byte_counter[1], n214) ;   // sha_top.v(226)
    assign sha_core_block_read_data_next[375] = n817 ? xram_data_in[7] : sha_core_block[375];   // sha_top.v(226)
    assign sha_core_block_read_data_next[374] = n817 ? xram_data_in[6] : sha_core_block[374];   // sha_top.v(226)
    assign sha_core_block_read_data_next[373] = n817 ? xram_data_in[5] : sha_core_block[373];   // sha_top.v(226)
    assign sha_core_block_read_data_next[372] = n817 ? xram_data_in[4] : sha_core_block[372];   // sha_top.v(226)
    assign sha_core_block_read_data_next[371] = n817 ? xram_data_in[3] : sha_core_block[371];   // sha_top.v(226)
    assign sha_core_block_read_data_next[370] = n817 ? xram_data_in[2] : sha_core_block[370];   // sha_top.v(226)
    assign sha_core_block_read_data_next[369] = n817 ? xram_data_in[1] : sha_core_block[369];   // sha_top.v(226)
    assign sha_core_block_read_data_next[368] = n817 ? xram_data_in[0] : sha_core_block[368];   // sha_top.v(226)
    nor (n827, byte_counter[5], n218, byte_counter[3], byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // sha_top.v(227)
    assign sha_core_block_read_data_next[383] = n827 ? xram_data_in[7] : sha_core_block[383];   // sha_top.v(227)
    assign sha_core_block_read_data_next[382] = n827 ? xram_data_in[6] : sha_core_block[382];   // sha_top.v(227)
    assign sha_core_block_read_data_next[381] = n827 ? xram_data_in[5] : sha_core_block[381];   // sha_top.v(227)
    assign sha_core_block_read_data_next[380] = n827 ? xram_data_in[4] : sha_core_block[380];   // sha_top.v(227)
    assign sha_core_block_read_data_next[379] = n827 ? xram_data_in[3] : sha_core_block[379];   // sha_top.v(227)
    assign sha_core_block_read_data_next[378] = n827 ? xram_data_in[2] : sha_core_block[378];   // sha_top.v(227)
    assign sha_core_block_read_data_next[377] = n827 ? xram_data_in[1] : sha_core_block[377];   // sha_top.v(227)
    assign sha_core_block_read_data_next[376] = n827 ? xram_data_in[0] : sha_core_block[376];   // sha_top.v(227)
    nor (n840, byte_counter[5], byte_counter[4], n217, n216, n215, 
        n214) ;   // sha_top.v(228)
    assign sha_core_block_read_data_next[391] = n840 ? xram_data_in[7] : sha_core_block[391];   // sha_top.v(228)
    assign sha_core_block_read_data_next[390] = n840 ? xram_data_in[6] : sha_core_block[390];   // sha_top.v(228)
    assign sha_core_block_read_data_next[389] = n840 ? xram_data_in[5] : sha_core_block[389];   // sha_top.v(228)
    assign sha_core_block_read_data_next[388] = n840 ? xram_data_in[4] : sha_core_block[388];   // sha_top.v(228)
    assign sha_core_block_read_data_next[387] = n840 ? xram_data_in[3] : sha_core_block[387];   // sha_top.v(228)
    assign sha_core_block_read_data_next[386] = n840 ? xram_data_in[2] : sha_core_block[386];   // sha_top.v(228)
    assign sha_core_block_read_data_next[385] = n840 ? xram_data_in[1] : sha_core_block[385];   // sha_top.v(228)
    assign sha_core_block_read_data_next[384] = n840 ? xram_data_in[0] : sha_core_block[384];   // sha_top.v(228)
    nor (n852, byte_counter[5], byte_counter[4], n217, n216, n215, 
        byte_counter[0]) ;   // sha_top.v(229)
    assign sha_core_block_read_data_next[399] = n852 ? xram_data_in[7] : sha_core_block[399];   // sha_top.v(229)
    assign sha_core_block_read_data_next[398] = n852 ? xram_data_in[6] : sha_core_block[398];   // sha_top.v(229)
    assign sha_core_block_read_data_next[397] = n852 ? xram_data_in[5] : sha_core_block[397];   // sha_top.v(229)
    assign sha_core_block_read_data_next[396] = n852 ? xram_data_in[4] : sha_core_block[396];   // sha_top.v(229)
    assign sha_core_block_read_data_next[395] = n852 ? xram_data_in[3] : sha_core_block[395];   // sha_top.v(229)
    assign sha_core_block_read_data_next[394] = n852 ? xram_data_in[2] : sha_core_block[394];   // sha_top.v(229)
    assign sha_core_block_read_data_next[393] = n852 ? xram_data_in[1] : sha_core_block[393];   // sha_top.v(229)
    assign sha_core_block_read_data_next[392] = n852 ? xram_data_in[0] : sha_core_block[392];   // sha_top.v(229)
    nor (n864, byte_counter[5], byte_counter[4], n217, n216, byte_counter[1], 
        n214) ;   // sha_top.v(230)
    assign sha_core_block_read_data_next[407] = n864 ? xram_data_in[7] : sha_core_block[407];   // sha_top.v(230)
    assign sha_core_block_read_data_next[406] = n864 ? xram_data_in[6] : sha_core_block[406];   // sha_top.v(230)
    assign sha_core_block_read_data_next[405] = n864 ? xram_data_in[5] : sha_core_block[405];   // sha_top.v(230)
    assign sha_core_block_read_data_next[404] = n864 ? xram_data_in[4] : sha_core_block[404];   // sha_top.v(230)
    assign sha_core_block_read_data_next[403] = n864 ? xram_data_in[3] : sha_core_block[403];   // sha_top.v(230)
    assign sha_core_block_read_data_next[402] = n864 ? xram_data_in[2] : sha_core_block[402];   // sha_top.v(230)
    assign sha_core_block_read_data_next[401] = n864 ? xram_data_in[1] : sha_core_block[401];   // sha_top.v(230)
    assign sha_core_block_read_data_next[400] = n864 ? xram_data_in[0] : sha_core_block[400];   // sha_top.v(230)
    nor (n875, byte_counter[5], byte_counter[4], n217, n216, byte_counter[1], 
        byte_counter[0]) ;   // sha_top.v(231)
    assign sha_core_block_read_data_next[415] = n875 ? xram_data_in[7] : sha_core_block[415];   // sha_top.v(231)
    assign sha_core_block_read_data_next[414] = n875 ? xram_data_in[6] : sha_core_block[414];   // sha_top.v(231)
    assign sha_core_block_read_data_next[413] = n875 ? xram_data_in[5] : sha_core_block[413];   // sha_top.v(231)
    assign sha_core_block_read_data_next[412] = n875 ? xram_data_in[4] : sha_core_block[412];   // sha_top.v(231)
    assign sha_core_block_read_data_next[411] = n875 ? xram_data_in[3] : sha_core_block[411];   // sha_top.v(231)
    assign sha_core_block_read_data_next[410] = n875 ? xram_data_in[2] : sha_core_block[410];   // sha_top.v(231)
    assign sha_core_block_read_data_next[409] = n875 ? xram_data_in[1] : sha_core_block[409];   // sha_top.v(231)
    assign sha_core_block_read_data_next[408] = n875 ? xram_data_in[0] : sha_core_block[408];   // sha_top.v(231)
    nor (n887, byte_counter[5], byte_counter[4], n217, byte_counter[2], 
        n215, n214) ;   // sha_top.v(232)
    assign sha_core_block_read_data_next[423] = n887 ? xram_data_in[7] : sha_core_block[423];   // sha_top.v(232)
    assign sha_core_block_read_data_next[422] = n887 ? xram_data_in[6] : sha_core_block[422];   // sha_top.v(232)
    assign sha_core_block_read_data_next[421] = n887 ? xram_data_in[5] : sha_core_block[421];   // sha_top.v(232)
    assign sha_core_block_read_data_next[420] = n887 ? xram_data_in[4] : sha_core_block[420];   // sha_top.v(232)
    assign sha_core_block_read_data_next[419] = n887 ? xram_data_in[3] : sha_core_block[419];   // sha_top.v(232)
    assign sha_core_block_read_data_next[418] = n887 ? xram_data_in[2] : sha_core_block[418];   // sha_top.v(232)
    assign sha_core_block_read_data_next[417] = n887 ? xram_data_in[1] : sha_core_block[417];   // sha_top.v(232)
    assign sha_core_block_read_data_next[416] = n887 ? xram_data_in[0] : sha_core_block[416];   // sha_top.v(232)
    nor (n898, byte_counter[5], byte_counter[4], n217, byte_counter[2], 
        n215, byte_counter[0]) ;   // sha_top.v(233)
    assign sha_core_block_read_data_next[431] = n898 ? xram_data_in[7] : sha_core_block[431];   // sha_top.v(233)
    assign sha_core_block_read_data_next[430] = n898 ? xram_data_in[6] : sha_core_block[430];   // sha_top.v(233)
    assign sha_core_block_read_data_next[429] = n898 ? xram_data_in[5] : sha_core_block[429];   // sha_top.v(233)
    assign sha_core_block_read_data_next[428] = n898 ? xram_data_in[4] : sha_core_block[428];   // sha_top.v(233)
    assign sha_core_block_read_data_next[427] = n898 ? xram_data_in[3] : sha_core_block[427];   // sha_top.v(233)
    assign sha_core_block_read_data_next[426] = n898 ? xram_data_in[2] : sha_core_block[426];   // sha_top.v(233)
    assign sha_core_block_read_data_next[425] = n898 ? xram_data_in[1] : sha_core_block[425];   // sha_top.v(233)
    assign sha_core_block_read_data_next[424] = n898 ? xram_data_in[0] : sha_core_block[424];   // sha_top.v(233)
    nor (n909, byte_counter[5], byte_counter[4], n217, byte_counter[2], 
        byte_counter[1], n214) ;   // sha_top.v(234)
    assign sha_core_block_read_data_next[439] = n909 ? xram_data_in[7] : sha_core_block[439];   // sha_top.v(234)
    assign sha_core_block_read_data_next[438] = n909 ? xram_data_in[6] : sha_core_block[438];   // sha_top.v(234)
    assign sha_core_block_read_data_next[437] = n909 ? xram_data_in[5] : sha_core_block[437];   // sha_top.v(234)
    assign sha_core_block_read_data_next[436] = n909 ? xram_data_in[4] : sha_core_block[436];   // sha_top.v(234)
    assign sha_core_block_read_data_next[435] = n909 ? xram_data_in[3] : sha_core_block[435];   // sha_top.v(234)
    assign sha_core_block_read_data_next[434] = n909 ? xram_data_in[2] : sha_core_block[434];   // sha_top.v(234)
    assign sha_core_block_read_data_next[433] = n909 ? xram_data_in[1] : sha_core_block[433];   // sha_top.v(234)
    assign sha_core_block_read_data_next[432] = n909 ? xram_data_in[0] : sha_core_block[432];   // sha_top.v(234)
    nor (n919, byte_counter[5], byte_counter[4], n217, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // sha_top.v(235)
    assign sha_core_block_read_data_next[447] = n919 ? xram_data_in[7] : sha_core_block[447];   // sha_top.v(235)
    assign sha_core_block_read_data_next[446] = n919 ? xram_data_in[6] : sha_core_block[446];   // sha_top.v(235)
    assign sha_core_block_read_data_next[445] = n919 ? xram_data_in[5] : sha_core_block[445];   // sha_top.v(235)
    assign sha_core_block_read_data_next[444] = n919 ? xram_data_in[4] : sha_core_block[444];   // sha_top.v(235)
    assign sha_core_block_read_data_next[443] = n919 ? xram_data_in[3] : sha_core_block[443];   // sha_top.v(235)
    assign sha_core_block_read_data_next[442] = n919 ? xram_data_in[2] : sha_core_block[442];   // sha_top.v(235)
    assign sha_core_block_read_data_next[441] = n919 ? xram_data_in[1] : sha_core_block[441];   // sha_top.v(235)
    assign sha_core_block_read_data_next[440] = n919 ? xram_data_in[0] : sha_core_block[440];   // sha_top.v(235)
    nor (n931, byte_counter[5], byte_counter[4], byte_counter[3], n216, 
        n215, n214) ;   // sha_top.v(236)
    assign sha_core_block_read_data_next[455] = n931 ? xram_data_in[7] : sha_core_block[455];   // sha_top.v(236)
    assign sha_core_block_read_data_next[454] = n931 ? xram_data_in[6] : sha_core_block[454];   // sha_top.v(236)
    assign sha_core_block_read_data_next[453] = n931 ? xram_data_in[5] : sha_core_block[453];   // sha_top.v(236)
    assign sha_core_block_read_data_next[452] = n931 ? xram_data_in[4] : sha_core_block[452];   // sha_top.v(236)
    assign sha_core_block_read_data_next[451] = n931 ? xram_data_in[3] : sha_core_block[451];   // sha_top.v(236)
    assign sha_core_block_read_data_next[450] = n931 ? xram_data_in[2] : sha_core_block[450];   // sha_top.v(236)
    assign sha_core_block_read_data_next[449] = n931 ? xram_data_in[1] : sha_core_block[449];   // sha_top.v(236)
    assign sha_core_block_read_data_next[448] = n931 ? xram_data_in[0] : sha_core_block[448];   // sha_top.v(236)
    nor (n942, byte_counter[5], byte_counter[4], byte_counter[3], n216, 
        n215, byte_counter[0]) ;   // sha_top.v(237)
    assign sha_core_block_read_data_next[463] = n942 ? xram_data_in[7] : sha_core_block[463];   // sha_top.v(237)
    assign sha_core_block_read_data_next[462] = n942 ? xram_data_in[6] : sha_core_block[462];   // sha_top.v(237)
    assign sha_core_block_read_data_next[461] = n942 ? xram_data_in[5] : sha_core_block[461];   // sha_top.v(237)
    assign sha_core_block_read_data_next[460] = n942 ? xram_data_in[4] : sha_core_block[460];   // sha_top.v(237)
    assign sha_core_block_read_data_next[459] = n942 ? xram_data_in[3] : sha_core_block[459];   // sha_top.v(237)
    assign sha_core_block_read_data_next[458] = n942 ? xram_data_in[2] : sha_core_block[458];   // sha_top.v(237)
    assign sha_core_block_read_data_next[457] = n942 ? xram_data_in[1] : sha_core_block[457];   // sha_top.v(237)
    assign sha_core_block_read_data_next[456] = n942 ? xram_data_in[0] : sha_core_block[456];   // sha_top.v(237)
    nor (n953, byte_counter[5], byte_counter[4], byte_counter[3], n216, 
        byte_counter[1], n214) ;   // sha_top.v(238)
    assign sha_core_block_read_data_next[471] = n953 ? xram_data_in[7] : sha_core_block[471];   // sha_top.v(238)
    assign sha_core_block_read_data_next[470] = n953 ? xram_data_in[6] : sha_core_block[470];   // sha_top.v(238)
    assign sha_core_block_read_data_next[469] = n953 ? xram_data_in[5] : sha_core_block[469];   // sha_top.v(238)
    assign sha_core_block_read_data_next[468] = n953 ? xram_data_in[4] : sha_core_block[468];   // sha_top.v(238)
    assign sha_core_block_read_data_next[467] = n953 ? xram_data_in[3] : sha_core_block[467];   // sha_top.v(238)
    assign sha_core_block_read_data_next[466] = n953 ? xram_data_in[2] : sha_core_block[466];   // sha_top.v(238)
    assign sha_core_block_read_data_next[465] = n953 ? xram_data_in[1] : sha_core_block[465];   // sha_top.v(238)
    assign sha_core_block_read_data_next[464] = n953 ? xram_data_in[0] : sha_core_block[464];   // sha_top.v(238)
    nor (n963, byte_counter[5], byte_counter[4], byte_counter[3], n216, 
        byte_counter[1], byte_counter[0]) ;   // sha_top.v(239)
    assign sha_core_block_read_data_next[479] = n963 ? xram_data_in[7] : sha_core_block[479];   // sha_top.v(239)
    assign sha_core_block_read_data_next[478] = n963 ? xram_data_in[6] : sha_core_block[478];   // sha_top.v(239)
    assign sha_core_block_read_data_next[477] = n963 ? xram_data_in[5] : sha_core_block[477];   // sha_top.v(239)
    assign sha_core_block_read_data_next[476] = n963 ? xram_data_in[4] : sha_core_block[476];   // sha_top.v(239)
    assign sha_core_block_read_data_next[475] = n963 ? xram_data_in[3] : sha_core_block[475];   // sha_top.v(239)
    assign sha_core_block_read_data_next[474] = n963 ? xram_data_in[2] : sha_core_block[474];   // sha_top.v(239)
    assign sha_core_block_read_data_next[473] = n963 ? xram_data_in[1] : sha_core_block[473];   // sha_top.v(239)
    assign sha_core_block_read_data_next[472] = n963 ? xram_data_in[0] : sha_core_block[472];   // sha_top.v(239)
    nor (n974, byte_counter[5], byte_counter[4], byte_counter[3], byte_counter[2], 
        n215, n214) ;   // sha_top.v(240)
    assign sha_core_block_read_data_next[487] = n974 ? xram_data_in[7] : sha_core_block[487];   // sha_top.v(240)
    assign sha_core_block_read_data_next[486] = n974 ? xram_data_in[6] : sha_core_block[486];   // sha_top.v(240)
    assign sha_core_block_read_data_next[485] = n974 ? xram_data_in[5] : sha_core_block[485];   // sha_top.v(240)
    assign sha_core_block_read_data_next[484] = n974 ? xram_data_in[4] : sha_core_block[484];   // sha_top.v(240)
    assign sha_core_block_read_data_next[483] = n974 ? xram_data_in[3] : sha_core_block[483];   // sha_top.v(240)
    assign sha_core_block_read_data_next[482] = n974 ? xram_data_in[2] : sha_core_block[482];   // sha_top.v(240)
    assign sha_core_block_read_data_next[481] = n974 ? xram_data_in[1] : sha_core_block[481];   // sha_top.v(240)
    assign sha_core_block_read_data_next[480] = n974 ? xram_data_in[0] : sha_core_block[480];   // sha_top.v(240)
    nor (n984, byte_counter[5], byte_counter[4], byte_counter[3], byte_counter[2], 
        n215, byte_counter[0]) ;   // sha_top.v(241)
    assign sha_core_block_read_data_next[495] = n984 ? xram_data_in[7] : sha_core_block[495];   // sha_top.v(241)
    assign sha_core_block_read_data_next[494] = n984 ? xram_data_in[6] : sha_core_block[494];   // sha_top.v(241)
    assign sha_core_block_read_data_next[493] = n984 ? xram_data_in[5] : sha_core_block[493];   // sha_top.v(241)
    assign sha_core_block_read_data_next[492] = n984 ? xram_data_in[4] : sha_core_block[492];   // sha_top.v(241)
    assign sha_core_block_read_data_next[491] = n984 ? xram_data_in[3] : sha_core_block[491];   // sha_top.v(241)
    assign sha_core_block_read_data_next[490] = n984 ? xram_data_in[2] : sha_core_block[490];   // sha_top.v(241)
    assign sha_core_block_read_data_next[489] = n984 ? xram_data_in[1] : sha_core_block[489];   // sha_top.v(241)
    assign sha_core_block_read_data_next[488] = n984 ? xram_data_in[0] : sha_core_block[488];   // sha_top.v(241)
    nor (n994, byte_counter[5], byte_counter[4], byte_counter[3], byte_counter[2], 
        byte_counter[1], n214) ;   // sha_top.v(242)
    assign sha_core_block_read_data_next[503] = n994 ? xram_data_in[7] : sha_core_block[503];   // sha_top.v(242)
    assign sha_core_block_read_data_next[502] = n994 ? xram_data_in[6] : sha_core_block[502];   // sha_top.v(242)
    assign sha_core_block_read_data_next[501] = n994 ? xram_data_in[5] : sha_core_block[501];   // sha_top.v(242)
    assign sha_core_block_read_data_next[500] = n994 ? xram_data_in[4] : sha_core_block[500];   // sha_top.v(242)
    assign sha_core_block_read_data_next[499] = n994 ? xram_data_in[3] : sha_core_block[499];   // sha_top.v(242)
    assign sha_core_block_read_data_next[498] = n994 ? xram_data_in[2] : sha_core_block[498];   // sha_top.v(242)
    assign sha_core_block_read_data_next[497] = n994 ? xram_data_in[1] : sha_core_block[497];   // sha_top.v(242)
    assign sha_core_block_read_data_next[496] = n994 ? xram_data_in[0] : sha_core_block[496];   // sha_top.v(242)
    nor (n1003, byte_counter[5], byte_counter[4], byte_counter[3], byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // sha_top.v(243)
    assign sha_core_block_read_data_next[511] = n1003 ? xram_data_in[7] : sha_core_block[511];   // sha_top.v(243)
    assign sha_core_block_read_data_next[510] = n1003 ? xram_data_in[6] : sha_core_block[510];   // sha_top.v(243)
    assign sha_core_block_read_data_next[509] = n1003 ? xram_data_in[5] : sha_core_block[509];   // sha_top.v(243)
    assign sha_core_block_read_data_next[508] = n1003 ? xram_data_in[4] : sha_core_block[508];   // sha_top.v(243)
    assign sha_core_block_read_data_next[507] = n1003 ? xram_data_in[3] : sha_core_block[507];   // sha_top.v(243)
    assign sha_core_block_read_data_next[506] = n1003 ? xram_data_in[2] : sha_core_block[506];   // sha_top.v(243)
    assign sha_core_block_read_data_next[505] = n1003 ? xram_data_in[1] : sha_core_block[505];   // sha_top.v(243)
    assign sha_core_block_read_data_next[504] = n1003 ? xram_data_in[0] : sha_core_block[504];   // sha_top.v(243)
    assign n1012 = sha_state_read_data ? sha_core_block_read_data_next[511] : sha_core_block[511];   // sha_top.v(246)
    assign n1013 = sha_state_read_data ? sha_core_block_read_data_next[510] : sha_core_block[510];   // sha_top.v(246)
    assign n1014 = sha_state_read_data ? sha_core_block_read_data_next[509] : sha_core_block[509];   // sha_top.v(246)
    assign n1015 = sha_state_read_data ? sha_core_block_read_data_next[508] : sha_core_block[508];   // sha_top.v(246)
    assign n1016 = sha_state_read_data ? sha_core_block_read_data_next[507] : sha_core_block[507];   // sha_top.v(246)
    assign n1017 = sha_state_read_data ? sha_core_block_read_data_next[506] : sha_core_block[506];   // sha_top.v(246)
    assign n1018 = sha_state_read_data ? sha_core_block_read_data_next[505] : sha_core_block[505];   // sha_top.v(246)
    assign n1019 = sha_state_read_data ? sha_core_block_read_data_next[504] : sha_core_block[504];   // sha_top.v(246)
    assign n1020 = sha_state_read_data ? sha_core_block_read_data_next[503] : sha_core_block[503];   // sha_top.v(246)
    assign n1021 = sha_state_read_data ? sha_core_block_read_data_next[502] : sha_core_block[502];   // sha_top.v(246)
    assign n1022 = sha_state_read_data ? sha_core_block_read_data_next[501] : sha_core_block[501];   // sha_top.v(246)
    assign n1023 = sha_state_read_data ? sha_core_block_read_data_next[500] : sha_core_block[500];   // sha_top.v(246)
    assign n1024 = sha_state_read_data ? sha_core_block_read_data_next[499] : sha_core_block[499];   // sha_top.v(246)
    assign n1025 = sha_state_read_data ? sha_core_block_read_data_next[498] : sha_core_block[498];   // sha_top.v(246)
    assign n1026 = sha_state_read_data ? sha_core_block_read_data_next[497] : sha_core_block[497];   // sha_top.v(246)
    assign n1027 = sha_state_read_data ? sha_core_block_read_data_next[496] : sha_core_block[496];   // sha_top.v(246)
    assign n1028 = sha_state_read_data ? sha_core_block_read_data_next[495] : sha_core_block[495];   // sha_top.v(246)
    assign n1029 = sha_state_read_data ? sha_core_block_read_data_next[494] : sha_core_block[494];   // sha_top.v(246)
    assign n1030 = sha_state_read_data ? sha_core_block_read_data_next[493] : sha_core_block[493];   // sha_top.v(246)
    assign n1031 = sha_state_read_data ? sha_core_block_read_data_next[492] : sha_core_block[492];   // sha_top.v(246)
    assign n1032 = sha_state_read_data ? sha_core_block_read_data_next[491] : sha_core_block[491];   // sha_top.v(246)
    assign n1033 = sha_state_read_data ? sha_core_block_read_data_next[490] : sha_core_block[490];   // sha_top.v(246)
    assign n1034 = sha_state_read_data ? sha_core_block_read_data_next[489] : sha_core_block[489];   // sha_top.v(246)
    assign n1035 = sha_state_read_data ? sha_core_block_read_data_next[488] : sha_core_block[488];   // sha_top.v(246)
    assign n1036 = sha_state_read_data ? sha_core_block_read_data_next[487] : sha_core_block[487];   // sha_top.v(246)
    assign n1037 = sha_state_read_data ? sha_core_block_read_data_next[486] : sha_core_block[486];   // sha_top.v(246)
    assign n1038 = sha_state_read_data ? sha_core_block_read_data_next[485] : sha_core_block[485];   // sha_top.v(246)
    assign n1039 = sha_state_read_data ? sha_core_block_read_data_next[484] : sha_core_block[484];   // sha_top.v(246)
    assign n1040 = sha_state_read_data ? sha_core_block_read_data_next[483] : sha_core_block[483];   // sha_top.v(246)
    assign n1041 = sha_state_read_data ? sha_core_block_read_data_next[482] : sha_core_block[482];   // sha_top.v(246)
    assign n1042 = sha_state_read_data ? sha_core_block_read_data_next[481] : sha_core_block[481];   // sha_top.v(246)
    assign n1043 = sha_state_read_data ? sha_core_block_read_data_next[480] : sha_core_block[480];   // sha_top.v(246)
    assign n1044 = sha_state_read_data ? sha_core_block_read_data_next[479] : sha_core_block[479];   // sha_top.v(246)
    assign n1045 = sha_state_read_data ? sha_core_block_read_data_next[478] : sha_core_block[478];   // sha_top.v(246)
    assign n1046 = sha_state_read_data ? sha_core_block_read_data_next[477] : sha_core_block[477];   // sha_top.v(246)
    assign n1047 = sha_state_read_data ? sha_core_block_read_data_next[476] : sha_core_block[476];   // sha_top.v(246)
    assign n1048 = sha_state_read_data ? sha_core_block_read_data_next[475] : sha_core_block[475];   // sha_top.v(246)
    assign n1049 = sha_state_read_data ? sha_core_block_read_data_next[474] : sha_core_block[474];   // sha_top.v(246)
    assign n1050 = sha_state_read_data ? sha_core_block_read_data_next[473] : sha_core_block[473];   // sha_top.v(246)
    assign n1051 = sha_state_read_data ? sha_core_block_read_data_next[472] : sha_core_block[472];   // sha_top.v(246)
    assign n1052 = sha_state_read_data ? sha_core_block_read_data_next[471] : sha_core_block[471];   // sha_top.v(246)
    assign n1053 = sha_state_read_data ? sha_core_block_read_data_next[470] : sha_core_block[470];   // sha_top.v(246)
    assign n1054 = sha_state_read_data ? sha_core_block_read_data_next[469] : sha_core_block[469];   // sha_top.v(246)
    assign n1055 = sha_state_read_data ? sha_core_block_read_data_next[468] : sha_core_block[468];   // sha_top.v(246)
    assign n1056 = sha_state_read_data ? sha_core_block_read_data_next[467] : sha_core_block[467];   // sha_top.v(246)
    assign n1057 = sha_state_read_data ? sha_core_block_read_data_next[466] : sha_core_block[466];   // sha_top.v(246)
    assign n1058 = sha_state_read_data ? sha_core_block_read_data_next[465] : sha_core_block[465];   // sha_top.v(246)
    assign n1059 = sha_state_read_data ? sha_core_block_read_data_next[464] : sha_core_block[464];   // sha_top.v(246)
    assign n1060 = sha_state_read_data ? sha_core_block_read_data_next[463] : sha_core_block[463];   // sha_top.v(246)
    assign n1061 = sha_state_read_data ? sha_core_block_read_data_next[462] : sha_core_block[462];   // sha_top.v(246)
    assign n1062 = sha_state_read_data ? sha_core_block_read_data_next[461] : sha_core_block[461];   // sha_top.v(246)
    assign n1063 = sha_state_read_data ? sha_core_block_read_data_next[460] : sha_core_block[460];   // sha_top.v(246)
    assign n1064 = sha_state_read_data ? sha_core_block_read_data_next[459] : sha_core_block[459];   // sha_top.v(246)
    assign n1065 = sha_state_read_data ? sha_core_block_read_data_next[458] : sha_core_block[458];   // sha_top.v(246)
    assign n1066 = sha_state_read_data ? sha_core_block_read_data_next[457] : sha_core_block[457];   // sha_top.v(246)
    assign n1067 = sha_state_read_data ? sha_core_block_read_data_next[456] : sha_core_block[456];   // sha_top.v(246)
    assign n1068 = sha_state_read_data ? sha_core_block_read_data_next[455] : sha_core_block[455];   // sha_top.v(246)
    assign n1069 = sha_state_read_data ? sha_core_block_read_data_next[454] : sha_core_block[454];   // sha_top.v(246)
    assign n1070 = sha_state_read_data ? sha_core_block_read_data_next[453] : sha_core_block[453];   // sha_top.v(246)
    assign n1071 = sha_state_read_data ? sha_core_block_read_data_next[452] : sha_core_block[452];   // sha_top.v(246)
    assign n1072 = sha_state_read_data ? sha_core_block_read_data_next[451] : sha_core_block[451];   // sha_top.v(246)
    assign n1073 = sha_state_read_data ? sha_core_block_read_data_next[450] : sha_core_block[450];   // sha_top.v(246)
    assign n1074 = sha_state_read_data ? sha_core_block_read_data_next[449] : sha_core_block[449];   // sha_top.v(246)
    assign n1075 = sha_state_read_data ? sha_core_block_read_data_next[448] : sha_core_block[448];   // sha_top.v(246)
    assign n1076 = sha_state_read_data ? sha_core_block_read_data_next[447] : sha_core_block[447];   // sha_top.v(246)
    assign n1077 = sha_state_read_data ? sha_core_block_read_data_next[446] : sha_core_block[446];   // sha_top.v(246)
    assign n1078 = sha_state_read_data ? sha_core_block_read_data_next[445] : sha_core_block[445];   // sha_top.v(246)
    assign n1079 = sha_state_read_data ? sha_core_block_read_data_next[444] : sha_core_block[444];   // sha_top.v(246)
    assign n1080 = sha_state_read_data ? sha_core_block_read_data_next[443] : sha_core_block[443];   // sha_top.v(246)
    assign n1081 = sha_state_read_data ? sha_core_block_read_data_next[442] : sha_core_block[442];   // sha_top.v(246)
    assign n1082 = sha_state_read_data ? sha_core_block_read_data_next[441] : sha_core_block[441];   // sha_top.v(246)
    assign n1083 = sha_state_read_data ? sha_core_block_read_data_next[440] : sha_core_block[440];   // sha_top.v(246)
    assign n1084 = sha_state_read_data ? sha_core_block_read_data_next[439] : sha_core_block[439];   // sha_top.v(246)
    assign n1085 = sha_state_read_data ? sha_core_block_read_data_next[438] : sha_core_block[438];   // sha_top.v(246)
    assign n1086 = sha_state_read_data ? sha_core_block_read_data_next[437] : sha_core_block[437];   // sha_top.v(246)
    assign n1087 = sha_state_read_data ? sha_core_block_read_data_next[436] : sha_core_block[436];   // sha_top.v(246)
    assign n1088 = sha_state_read_data ? sha_core_block_read_data_next[435] : sha_core_block[435];   // sha_top.v(246)
    assign n1089 = sha_state_read_data ? sha_core_block_read_data_next[434] : sha_core_block[434];   // sha_top.v(246)
    assign n1090 = sha_state_read_data ? sha_core_block_read_data_next[433] : sha_core_block[433];   // sha_top.v(246)
    assign n1091 = sha_state_read_data ? sha_core_block_read_data_next[432] : sha_core_block[432];   // sha_top.v(246)
    assign n1092 = sha_state_read_data ? sha_core_block_read_data_next[431] : sha_core_block[431];   // sha_top.v(246)
    assign n1093 = sha_state_read_data ? sha_core_block_read_data_next[430] : sha_core_block[430];   // sha_top.v(246)
    assign n1094 = sha_state_read_data ? sha_core_block_read_data_next[429] : sha_core_block[429];   // sha_top.v(246)
    assign n1095 = sha_state_read_data ? sha_core_block_read_data_next[428] : sha_core_block[428];   // sha_top.v(246)
    assign n1096 = sha_state_read_data ? sha_core_block_read_data_next[427] : sha_core_block[427];   // sha_top.v(246)
    assign n1097 = sha_state_read_data ? sha_core_block_read_data_next[426] : sha_core_block[426];   // sha_top.v(246)
    assign n1098 = sha_state_read_data ? sha_core_block_read_data_next[425] : sha_core_block[425];   // sha_top.v(246)
    assign n1099 = sha_state_read_data ? sha_core_block_read_data_next[424] : sha_core_block[424];   // sha_top.v(246)
    assign n1100 = sha_state_read_data ? sha_core_block_read_data_next[423] : sha_core_block[423];   // sha_top.v(246)
    assign n1101 = sha_state_read_data ? sha_core_block_read_data_next[422] : sha_core_block[422];   // sha_top.v(246)
    assign n1102 = sha_state_read_data ? sha_core_block_read_data_next[421] : sha_core_block[421];   // sha_top.v(246)
    assign n1103 = sha_state_read_data ? sha_core_block_read_data_next[420] : sha_core_block[420];   // sha_top.v(246)
    assign n1104 = sha_state_read_data ? sha_core_block_read_data_next[419] : sha_core_block[419];   // sha_top.v(246)
    assign n1105 = sha_state_read_data ? sha_core_block_read_data_next[418] : sha_core_block[418];   // sha_top.v(246)
    assign n1106 = sha_state_read_data ? sha_core_block_read_data_next[417] : sha_core_block[417];   // sha_top.v(246)
    assign n1107 = sha_state_read_data ? sha_core_block_read_data_next[416] : sha_core_block[416];   // sha_top.v(246)
    assign n1108 = sha_state_read_data ? sha_core_block_read_data_next[415] : sha_core_block[415];   // sha_top.v(246)
    assign n1109 = sha_state_read_data ? sha_core_block_read_data_next[414] : sha_core_block[414];   // sha_top.v(246)
    assign n1110 = sha_state_read_data ? sha_core_block_read_data_next[413] : sha_core_block[413];   // sha_top.v(246)
    assign n1111 = sha_state_read_data ? sha_core_block_read_data_next[412] : sha_core_block[412];   // sha_top.v(246)
    assign n1112 = sha_state_read_data ? sha_core_block_read_data_next[411] : sha_core_block[411];   // sha_top.v(246)
    assign n1113 = sha_state_read_data ? sha_core_block_read_data_next[410] : sha_core_block[410];   // sha_top.v(246)
    assign n1114 = sha_state_read_data ? sha_core_block_read_data_next[409] : sha_core_block[409];   // sha_top.v(246)
    assign n1115 = sha_state_read_data ? sha_core_block_read_data_next[408] : sha_core_block[408];   // sha_top.v(246)
    assign n1116 = sha_state_read_data ? sha_core_block_read_data_next[407] : sha_core_block[407];   // sha_top.v(246)
    assign n1117 = sha_state_read_data ? sha_core_block_read_data_next[406] : sha_core_block[406];   // sha_top.v(246)
    assign n1118 = sha_state_read_data ? sha_core_block_read_data_next[405] : sha_core_block[405];   // sha_top.v(246)
    assign n1119 = sha_state_read_data ? sha_core_block_read_data_next[404] : sha_core_block[404];   // sha_top.v(246)
    assign n1120 = sha_state_read_data ? sha_core_block_read_data_next[403] : sha_core_block[403];   // sha_top.v(246)
    assign n1121 = sha_state_read_data ? sha_core_block_read_data_next[402] : sha_core_block[402];   // sha_top.v(246)
    assign n1122 = sha_state_read_data ? sha_core_block_read_data_next[401] : sha_core_block[401];   // sha_top.v(246)
    assign n1123 = sha_state_read_data ? sha_core_block_read_data_next[400] : sha_core_block[400];   // sha_top.v(246)
    assign n1124 = sha_state_read_data ? sha_core_block_read_data_next[399] : sha_core_block[399];   // sha_top.v(246)
    assign n1125 = sha_state_read_data ? sha_core_block_read_data_next[398] : sha_core_block[398];   // sha_top.v(246)
    assign n1126 = sha_state_read_data ? sha_core_block_read_data_next[397] : sha_core_block[397];   // sha_top.v(246)
    assign n1127 = sha_state_read_data ? sha_core_block_read_data_next[396] : sha_core_block[396];   // sha_top.v(246)
    assign n1128 = sha_state_read_data ? sha_core_block_read_data_next[395] : sha_core_block[395];   // sha_top.v(246)
    assign n1129 = sha_state_read_data ? sha_core_block_read_data_next[394] : sha_core_block[394];   // sha_top.v(246)
    assign n1130 = sha_state_read_data ? sha_core_block_read_data_next[393] : sha_core_block[393];   // sha_top.v(246)
    assign n1131 = sha_state_read_data ? sha_core_block_read_data_next[392] : sha_core_block[392];   // sha_top.v(246)
    assign n1132 = sha_state_read_data ? sha_core_block_read_data_next[391] : sha_core_block[391];   // sha_top.v(246)
    assign n1133 = sha_state_read_data ? sha_core_block_read_data_next[390] : sha_core_block[390];   // sha_top.v(246)
    assign n1134 = sha_state_read_data ? sha_core_block_read_data_next[389] : sha_core_block[389];   // sha_top.v(246)
    assign n1135 = sha_state_read_data ? sha_core_block_read_data_next[388] : sha_core_block[388];   // sha_top.v(246)
    assign n1136 = sha_state_read_data ? sha_core_block_read_data_next[387] : sha_core_block[387];   // sha_top.v(246)
    assign n1137 = sha_state_read_data ? sha_core_block_read_data_next[386] : sha_core_block[386];   // sha_top.v(246)
    assign n1138 = sha_state_read_data ? sha_core_block_read_data_next[385] : sha_core_block[385];   // sha_top.v(246)
    assign n1139 = sha_state_read_data ? sha_core_block_read_data_next[384] : sha_core_block[384];   // sha_top.v(246)
    assign n1140 = sha_state_read_data ? sha_core_block_read_data_next[383] : sha_core_block[383];   // sha_top.v(246)
    assign n1141 = sha_state_read_data ? sha_core_block_read_data_next[382] : sha_core_block[382];   // sha_top.v(246)
    assign n1142 = sha_state_read_data ? sha_core_block_read_data_next[381] : sha_core_block[381];   // sha_top.v(246)
    assign n1143 = sha_state_read_data ? sha_core_block_read_data_next[380] : sha_core_block[380];   // sha_top.v(246)
    assign n1144 = sha_state_read_data ? sha_core_block_read_data_next[379] : sha_core_block[379];   // sha_top.v(246)
    assign n1145 = sha_state_read_data ? sha_core_block_read_data_next[378] : sha_core_block[378];   // sha_top.v(246)
    assign n1146 = sha_state_read_data ? sha_core_block_read_data_next[377] : sha_core_block[377];   // sha_top.v(246)
    assign n1147 = sha_state_read_data ? sha_core_block_read_data_next[376] : sha_core_block[376];   // sha_top.v(246)
    assign n1148 = sha_state_read_data ? sha_core_block_read_data_next[375] : sha_core_block[375];   // sha_top.v(246)
    assign n1149 = sha_state_read_data ? sha_core_block_read_data_next[374] : sha_core_block[374];   // sha_top.v(246)
    assign n1150 = sha_state_read_data ? sha_core_block_read_data_next[373] : sha_core_block[373];   // sha_top.v(246)
    assign n1151 = sha_state_read_data ? sha_core_block_read_data_next[372] : sha_core_block[372];   // sha_top.v(246)
    assign n1152 = sha_state_read_data ? sha_core_block_read_data_next[371] : sha_core_block[371];   // sha_top.v(246)
    assign n1153 = sha_state_read_data ? sha_core_block_read_data_next[370] : sha_core_block[370];   // sha_top.v(246)
    assign n1154 = sha_state_read_data ? sha_core_block_read_data_next[369] : sha_core_block[369];   // sha_top.v(246)
    assign n1155 = sha_state_read_data ? sha_core_block_read_data_next[368] : sha_core_block[368];   // sha_top.v(246)
    assign n1156 = sha_state_read_data ? sha_core_block_read_data_next[367] : sha_core_block[367];   // sha_top.v(246)
    assign n1157 = sha_state_read_data ? sha_core_block_read_data_next[366] : sha_core_block[366];   // sha_top.v(246)
    assign n1158 = sha_state_read_data ? sha_core_block_read_data_next[365] : sha_core_block[365];   // sha_top.v(246)
    assign n1159 = sha_state_read_data ? sha_core_block_read_data_next[364] : sha_core_block[364];   // sha_top.v(246)
    assign n1160 = sha_state_read_data ? sha_core_block_read_data_next[363] : sha_core_block[363];   // sha_top.v(246)
    assign n1161 = sha_state_read_data ? sha_core_block_read_data_next[362] : sha_core_block[362];   // sha_top.v(246)
    assign n1162 = sha_state_read_data ? sha_core_block_read_data_next[361] : sha_core_block[361];   // sha_top.v(246)
    assign n1163 = sha_state_read_data ? sha_core_block_read_data_next[360] : sha_core_block[360];   // sha_top.v(246)
    assign n1164 = sha_state_read_data ? sha_core_block_read_data_next[359] : sha_core_block[359];   // sha_top.v(246)
    assign n1165 = sha_state_read_data ? sha_core_block_read_data_next[358] : sha_core_block[358];   // sha_top.v(246)
    assign n1166 = sha_state_read_data ? sha_core_block_read_data_next[357] : sha_core_block[357];   // sha_top.v(246)
    assign n1167 = sha_state_read_data ? sha_core_block_read_data_next[356] : sha_core_block[356];   // sha_top.v(246)
    assign n1168 = sha_state_read_data ? sha_core_block_read_data_next[355] : sha_core_block[355];   // sha_top.v(246)
    assign n1169 = sha_state_read_data ? sha_core_block_read_data_next[354] : sha_core_block[354];   // sha_top.v(246)
    assign n1170 = sha_state_read_data ? sha_core_block_read_data_next[353] : sha_core_block[353];   // sha_top.v(246)
    assign n1171 = sha_state_read_data ? sha_core_block_read_data_next[352] : sha_core_block[352];   // sha_top.v(246)
    assign n1172 = sha_state_read_data ? sha_core_block_read_data_next[351] : sha_core_block[351];   // sha_top.v(246)
    assign n1173 = sha_state_read_data ? sha_core_block_read_data_next[350] : sha_core_block[350];   // sha_top.v(246)
    assign n1174 = sha_state_read_data ? sha_core_block_read_data_next[349] : sha_core_block[349];   // sha_top.v(246)
    assign n1175 = sha_state_read_data ? sha_core_block_read_data_next[348] : sha_core_block[348];   // sha_top.v(246)
    assign n1176 = sha_state_read_data ? sha_core_block_read_data_next[347] : sha_core_block[347];   // sha_top.v(246)
    assign n1177 = sha_state_read_data ? sha_core_block_read_data_next[346] : sha_core_block[346];   // sha_top.v(246)
    assign n1178 = sha_state_read_data ? sha_core_block_read_data_next[345] : sha_core_block[345];   // sha_top.v(246)
    assign n1179 = sha_state_read_data ? sha_core_block_read_data_next[344] : sha_core_block[344];   // sha_top.v(246)
    assign n1180 = sha_state_read_data ? sha_core_block_read_data_next[343] : sha_core_block[343];   // sha_top.v(246)
    assign n1181 = sha_state_read_data ? sha_core_block_read_data_next[342] : sha_core_block[342];   // sha_top.v(246)
    assign n1182 = sha_state_read_data ? sha_core_block_read_data_next[341] : sha_core_block[341];   // sha_top.v(246)
    assign n1183 = sha_state_read_data ? sha_core_block_read_data_next[340] : sha_core_block[340];   // sha_top.v(246)
    assign n1184 = sha_state_read_data ? sha_core_block_read_data_next[339] : sha_core_block[339];   // sha_top.v(246)
    assign n1185 = sha_state_read_data ? sha_core_block_read_data_next[338] : sha_core_block[338];   // sha_top.v(246)
    assign n1186 = sha_state_read_data ? sha_core_block_read_data_next[337] : sha_core_block[337];   // sha_top.v(246)
    assign n1187 = sha_state_read_data ? sha_core_block_read_data_next[336] : sha_core_block[336];   // sha_top.v(246)
    assign n1188 = sha_state_read_data ? sha_core_block_read_data_next[335] : sha_core_block[335];   // sha_top.v(246)
    assign n1189 = sha_state_read_data ? sha_core_block_read_data_next[334] : sha_core_block[334];   // sha_top.v(246)
    assign n1190 = sha_state_read_data ? sha_core_block_read_data_next[333] : sha_core_block[333];   // sha_top.v(246)
    assign n1191 = sha_state_read_data ? sha_core_block_read_data_next[332] : sha_core_block[332];   // sha_top.v(246)
    assign n1192 = sha_state_read_data ? sha_core_block_read_data_next[331] : sha_core_block[331];   // sha_top.v(246)
    assign n1193 = sha_state_read_data ? sha_core_block_read_data_next[330] : sha_core_block[330];   // sha_top.v(246)
    assign n1194 = sha_state_read_data ? sha_core_block_read_data_next[329] : sha_core_block[329];   // sha_top.v(246)
    assign n1195 = sha_state_read_data ? sha_core_block_read_data_next[328] : sha_core_block[328];   // sha_top.v(246)
    assign n1196 = sha_state_read_data ? sha_core_block_read_data_next[327] : sha_core_block[327];   // sha_top.v(246)
    assign n1197 = sha_state_read_data ? sha_core_block_read_data_next[326] : sha_core_block[326];   // sha_top.v(246)
    assign n1198 = sha_state_read_data ? sha_core_block_read_data_next[325] : sha_core_block[325];   // sha_top.v(246)
    assign n1199 = sha_state_read_data ? sha_core_block_read_data_next[324] : sha_core_block[324];   // sha_top.v(246)
    assign n1200 = sha_state_read_data ? sha_core_block_read_data_next[323] : sha_core_block[323];   // sha_top.v(246)
    assign n1201 = sha_state_read_data ? sha_core_block_read_data_next[322] : sha_core_block[322];   // sha_top.v(246)
    assign n1202 = sha_state_read_data ? sha_core_block_read_data_next[321] : sha_core_block[321];   // sha_top.v(246)
    assign n1203 = sha_state_read_data ? sha_core_block_read_data_next[320] : sha_core_block[320];   // sha_top.v(246)
    assign n1204 = sha_state_read_data ? sha_core_block_read_data_next[319] : sha_core_block[319];   // sha_top.v(246)
    assign n1205 = sha_state_read_data ? sha_core_block_read_data_next[318] : sha_core_block[318];   // sha_top.v(246)
    assign n1206 = sha_state_read_data ? sha_core_block_read_data_next[317] : sha_core_block[317];   // sha_top.v(246)
    assign n1207 = sha_state_read_data ? sha_core_block_read_data_next[316] : sha_core_block[316];   // sha_top.v(246)
    assign n1208 = sha_state_read_data ? sha_core_block_read_data_next[315] : sha_core_block[315];   // sha_top.v(246)
    assign n1209 = sha_state_read_data ? sha_core_block_read_data_next[314] : sha_core_block[314];   // sha_top.v(246)
    assign n1210 = sha_state_read_data ? sha_core_block_read_data_next[313] : sha_core_block[313];   // sha_top.v(246)
    assign n1211 = sha_state_read_data ? sha_core_block_read_data_next[312] : sha_core_block[312];   // sha_top.v(246)
    assign n1212 = sha_state_read_data ? sha_core_block_read_data_next[311] : sha_core_block[311];   // sha_top.v(246)
    assign n1213 = sha_state_read_data ? sha_core_block_read_data_next[310] : sha_core_block[310];   // sha_top.v(246)
    assign n1214 = sha_state_read_data ? sha_core_block_read_data_next[309] : sha_core_block[309];   // sha_top.v(246)
    assign n1215 = sha_state_read_data ? sha_core_block_read_data_next[308] : sha_core_block[308];   // sha_top.v(246)
    assign n1216 = sha_state_read_data ? sha_core_block_read_data_next[307] : sha_core_block[307];   // sha_top.v(246)
    assign n1217 = sha_state_read_data ? sha_core_block_read_data_next[306] : sha_core_block[306];   // sha_top.v(246)
    assign n1218 = sha_state_read_data ? sha_core_block_read_data_next[305] : sha_core_block[305];   // sha_top.v(246)
    assign n1219 = sha_state_read_data ? sha_core_block_read_data_next[304] : sha_core_block[304];   // sha_top.v(246)
    assign n1220 = sha_state_read_data ? sha_core_block_read_data_next[303] : sha_core_block[303];   // sha_top.v(246)
    assign n1221 = sha_state_read_data ? sha_core_block_read_data_next[302] : sha_core_block[302];   // sha_top.v(246)
    assign n1222 = sha_state_read_data ? sha_core_block_read_data_next[301] : sha_core_block[301];   // sha_top.v(246)
    assign n1223 = sha_state_read_data ? sha_core_block_read_data_next[300] : sha_core_block[300];   // sha_top.v(246)
    assign n1224 = sha_state_read_data ? sha_core_block_read_data_next[299] : sha_core_block[299];   // sha_top.v(246)
    assign n1225 = sha_state_read_data ? sha_core_block_read_data_next[298] : sha_core_block[298];   // sha_top.v(246)
    assign n1226 = sha_state_read_data ? sha_core_block_read_data_next[297] : sha_core_block[297];   // sha_top.v(246)
    assign n1227 = sha_state_read_data ? sha_core_block_read_data_next[296] : sha_core_block[296];   // sha_top.v(246)
    assign n1228 = sha_state_read_data ? sha_core_block_read_data_next[295] : sha_core_block[295];   // sha_top.v(246)
    assign n1229 = sha_state_read_data ? sha_core_block_read_data_next[294] : sha_core_block[294];   // sha_top.v(246)
    assign n1230 = sha_state_read_data ? sha_core_block_read_data_next[293] : sha_core_block[293];   // sha_top.v(246)
    assign n1231 = sha_state_read_data ? sha_core_block_read_data_next[292] : sha_core_block[292];   // sha_top.v(246)
    assign n1232 = sha_state_read_data ? sha_core_block_read_data_next[291] : sha_core_block[291];   // sha_top.v(246)
    assign n1233 = sha_state_read_data ? sha_core_block_read_data_next[290] : sha_core_block[290];   // sha_top.v(246)
    assign n1234 = sha_state_read_data ? sha_core_block_read_data_next[289] : sha_core_block[289];   // sha_top.v(246)
    assign n1235 = sha_state_read_data ? sha_core_block_read_data_next[288] : sha_core_block[288];   // sha_top.v(246)
    assign n1236 = sha_state_read_data ? sha_core_block_read_data_next[287] : sha_core_block[287];   // sha_top.v(246)
    assign n1237 = sha_state_read_data ? sha_core_block_read_data_next[286] : sha_core_block[286];   // sha_top.v(246)
    assign n1238 = sha_state_read_data ? sha_core_block_read_data_next[285] : sha_core_block[285];   // sha_top.v(246)
    assign n1239 = sha_state_read_data ? sha_core_block_read_data_next[284] : sha_core_block[284];   // sha_top.v(246)
    assign n1240 = sha_state_read_data ? sha_core_block_read_data_next[283] : sha_core_block[283];   // sha_top.v(246)
    assign n1241 = sha_state_read_data ? sha_core_block_read_data_next[282] : sha_core_block[282];   // sha_top.v(246)
    assign n1242 = sha_state_read_data ? sha_core_block_read_data_next[281] : sha_core_block[281];   // sha_top.v(246)
    assign n1243 = sha_state_read_data ? sha_core_block_read_data_next[280] : sha_core_block[280];   // sha_top.v(246)
    assign n1244 = sha_state_read_data ? sha_core_block_read_data_next[279] : sha_core_block[279];   // sha_top.v(246)
    assign n1245 = sha_state_read_data ? sha_core_block_read_data_next[278] : sha_core_block[278];   // sha_top.v(246)
    assign n1246 = sha_state_read_data ? sha_core_block_read_data_next[277] : sha_core_block[277];   // sha_top.v(246)
    assign n1247 = sha_state_read_data ? sha_core_block_read_data_next[276] : sha_core_block[276];   // sha_top.v(246)
    assign n1248 = sha_state_read_data ? sha_core_block_read_data_next[275] : sha_core_block[275];   // sha_top.v(246)
    assign n1249 = sha_state_read_data ? sha_core_block_read_data_next[274] : sha_core_block[274];   // sha_top.v(246)
    assign n1250 = sha_state_read_data ? sha_core_block_read_data_next[273] : sha_core_block[273];   // sha_top.v(246)
    assign n1251 = sha_state_read_data ? sha_core_block_read_data_next[272] : sha_core_block[272];   // sha_top.v(246)
    assign n1252 = sha_state_read_data ? sha_core_block_read_data_next[271] : sha_core_block[271];   // sha_top.v(246)
    assign n1253 = sha_state_read_data ? sha_core_block_read_data_next[270] : sha_core_block[270];   // sha_top.v(246)
    assign n1254 = sha_state_read_data ? sha_core_block_read_data_next[269] : sha_core_block[269];   // sha_top.v(246)
    assign n1255 = sha_state_read_data ? sha_core_block_read_data_next[268] : sha_core_block[268];   // sha_top.v(246)
    assign n1256 = sha_state_read_data ? sha_core_block_read_data_next[267] : sha_core_block[267];   // sha_top.v(246)
    assign n1257 = sha_state_read_data ? sha_core_block_read_data_next[266] : sha_core_block[266];   // sha_top.v(246)
    assign n1258 = sha_state_read_data ? sha_core_block_read_data_next[265] : sha_core_block[265];   // sha_top.v(246)
    assign n1259 = sha_state_read_data ? sha_core_block_read_data_next[264] : sha_core_block[264];   // sha_top.v(246)
    assign n1260 = sha_state_read_data ? sha_core_block_read_data_next[263] : sha_core_block[263];   // sha_top.v(246)
    assign n1261 = sha_state_read_data ? sha_core_block_read_data_next[262] : sha_core_block[262];   // sha_top.v(246)
    assign n1262 = sha_state_read_data ? sha_core_block_read_data_next[261] : sha_core_block[261];   // sha_top.v(246)
    assign n1263 = sha_state_read_data ? sha_core_block_read_data_next[260] : sha_core_block[260];   // sha_top.v(246)
    assign n1264 = sha_state_read_data ? sha_core_block_read_data_next[259] : sha_core_block[259];   // sha_top.v(246)
    assign n1265 = sha_state_read_data ? sha_core_block_read_data_next[258] : sha_core_block[258];   // sha_top.v(246)
    assign n1266 = sha_state_read_data ? sha_core_block_read_data_next[257] : sha_core_block[257];   // sha_top.v(246)
    assign n1267 = sha_state_read_data ? sha_core_block_read_data_next[256] : sha_core_block[256];   // sha_top.v(246)
    assign n1268 = sha_state_read_data ? sha_core_block_read_data_next[255] : sha_core_block[255];   // sha_top.v(246)
    assign n1269 = sha_state_read_data ? sha_core_block_read_data_next[254] : sha_core_block[254];   // sha_top.v(246)
    assign n1270 = sha_state_read_data ? sha_core_block_read_data_next[253] : sha_core_block[253];   // sha_top.v(246)
    assign n1271 = sha_state_read_data ? sha_core_block_read_data_next[252] : sha_core_block[252];   // sha_top.v(246)
    assign n1272 = sha_state_read_data ? sha_core_block_read_data_next[251] : sha_core_block[251];   // sha_top.v(246)
    assign n1273 = sha_state_read_data ? sha_core_block_read_data_next[250] : sha_core_block[250];   // sha_top.v(246)
    assign n1274 = sha_state_read_data ? sha_core_block_read_data_next[249] : sha_core_block[249];   // sha_top.v(246)
    assign n1275 = sha_state_read_data ? sha_core_block_read_data_next[248] : sha_core_block[248];   // sha_top.v(246)
    assign n1276 = sha_state_read_data ? sha_core_block_read_data_next[247] : sha_core_block[247];   // sha_top.v(246)
    assign n1277 = sha_state_read_data ? sha_core_block_read_data_next[246] : sha_core_block[246];   // sha_top.v(246)
    assign n1278 = sha_state_read_data ? sha_core_block_read_data_next[245] : sha_core_block[245];   // sha_top.v(246)
    assign n1279 = sha_state_read_data ? sha_core_block_read_data_next[244] : sha_core_block[244];   // sha_top.v(246)
    assign n1280 = sha_state_read_data ? sha_core_block_read_data_next[243] : sha_core_block[243];   // sha_top.v(246)
    assign n1281 = sha_state_read_data ? sha_core_block_read_data_next[242] : sha_core_block[242];   // sha_top.v(246)
    assign n1282 = sha_state_read_data ? sha_core_block_read_data_next[241] : sha_core_block[241];   // sha_top.v(246)
    assign n1283 = sha_state_read_data ? sha_core_block_read_data_next[240] : sha_core_block[240];   // sha_top.v(246)
    assign n1284 = sha_state_read_data ? sha_core_block_read_data_next[239] : sha_core_block[239];   // sha_top.v(246)
    assign n1285 = sha_state_read_data ? sha_core_block_read_data_next[238] : sha_core_block[238];   // sha_top.v(246)
    assign n1286 = sha_state_read_data ? sha_core_block_read_data_next[237] : sha_core_block[237];   // sha_top.v(246)
    assign n1287 = sha_state_read_data ? sha_core_block_read_data_next[236] : sha_core_block[236];   // sha_top.v(246)
    assign n1288 = sha_state_read_data ? sha_core_block_read_data_next[235] : sha_core_block[235];   // sha_top.v(246)
    assign n1289 = sha_state_read_data ? sha_core_block_read_data_next[234] : sha_core_block[234];   // sha_top.v(246)
    assign n1290 = sha_state_read_data ? sha_core_block_read_data_next[233] : sha_core_block[233];   // sha_top.v(246)
    assign n1291 = sha_state_read_data ? sha_core_block_read_data_next[232] : sha_core_block[232];   // sha_top.v(246)
    assign n1292 = sha_state_read_data ? sha_core_block_read_data_next[231] : sha_core_block[231];   // sha_top.v(246)
    assign n1293 = sha_state_read_data ? sha_core_block_read_data_next[230] : sha_core_block[230];   // sha_top.v(246)
    assign n1294 = sha_state_read_data ? sha_core_block_read_data_next[229] : sha_core_block[229];   // sha_top.v(246)
    assign n1295 = sha_state_read_data ? sha_core_block_read_data_next[228] : sha_core_block[228];   // sha_top.v(246)
    assign n1296 = sha_state_read_data ? sha_core_block_read_data_next[227] : sha_core_block[227];   // sha_top.v(246)
    assign n1297 = sha_state_read_data ? sha_core_block_read_data_next[226] : sha_core_block[226];   // sha_top.v(246)
    assign n1298 = sha_state_read_data ? sha_core_block_read_data_next[225] : sha_core_block[225];   // sha_top.v(246)
    assign n1299 = sha_state_read_data ? sha_core_block_read_data_next[224] : sha_core_block[224];   // sha_top.v(246)
    assign n1300 = sha_state_read_data ? sha_core_block_read_data_next[223] : sha_core_block[223];   // sha_top.v(246)
    assign n1301 = sha_state_read_data ? sha_core_block_read_data_next[222] : sha_core_block[222];   // sha_top.v(246)
    assign n1302 = sha_state_read_data ? sha_core_block_read_data_next[221] : sha_core_block[221];   // sha_top.v(246)
    assign n1303 = sha_state_read_data ? sha_core_block_read_data_next[220] : sha_core_block[220];   // sha_top.v(246)
    assign n1304 = sha_state_read_data ? sha_core_block_read_data_next[219] : sha_core_block[219];   // sha_top.v(246)
    assign n1305 = sha_state_read_data ? sha_core_block_read_data_next[218] : sha_core_block[218];   // sha_top.v(246)
    assign n1306 = sha_state_read_data ? sha_core_block_read_data_next[217] : sha_core_block[217];   // sha_top.v(246)
    assign n1307 = sha_state_read_data ? sha_core_block_read_data_next[216] : sha_core_block[216];   // sha_top.v(246)
    assign n1308 = sha_state_read_data ? sha_core_block_read_data_next[215] : sha_core_block[215];   // sha_top.v(246)
    assign n1309 = sha_state_read_data ? sha_core_block_read_data_next[214] : sha_core_block[214];   // sha_top.v(246)
    assign n1310 = sha_state_read_data ? sha_core_block_read_data_next[213] : sha_core_block[213];   // sha_top.v(246)
    assign n1311 = sha_state_read_data ? sha_core_block_read_data_next[212] : sha_core_block[212];   // sha_top.v(246)
    assign n1312 = sha_state_read_data ? sha_core_block_read_data_next[211] : sha_core_block[211];   // sha_top.v(246)
    assign n1313 = sha_state_read_data ? sha_core_block_read_data_next[210] : sha_core_block[210];   // sha_top.v(246)
    assign n1314 = sha_state_read_data ? sha_core_block_read_data_next[209] : sha_core_block[209];   // sha_top.v(246)
    assign n1315 = sha_state_read_data ? sha_core_block_read_data_next[208] : sha_core_block[208];   // sha_top.v(246)
    assign n1316 = sha_state_read_data ? sha_core_block_read_data_next[207] : sha_core_block[207];   // sha_top.v(246)
    assign n1317 = sha_state_read_data ? sha_core_block_read_data_next[206] : sha_core_block[206];   // sha_top.v(246)
    assign n1318 = sha_state_read_data ? sha_core_block_read_data_next[205] : sha_core_block[205];   // sha_top.v(246)
    assign n1319 = sha_state_read_data ? sha_core_block_read_data_next[204] : sha_core_block[204];   // sha_top.v(246)
    assign n1320 = sha_state_read_data ? sha_core_block_read_data_next[203] : sha_core_block[203];   // sha_top.v(246)
    assign n1321 = sha_state_read_data ? sha_core_block_read_data_next[202] : sha_core_block[202];   // sha_top.v(246)
    assign n1322 = sha_state_read_data ? sha_core_block_read_data_next[201] : sha_core_block[201];   // sha_top.v(246)
    assign n1323 = sha_state_read_data ? sha_core_block_read_data_next[200] : sha_core_block[200];   // sha_top.v(246)
    assign n1324 = sha_state_read_data ? sha_core_block_read_data_next[199] : sha_core_block[199];   // sha_top.v(246)
    assign n1325 = sha_state_read_data ? sha_core_block_read_data_next[198] : sha_core_block[198];   // sha_top.v(246)
    assign n1326 = sha_state_read_data ? sha_core_block_read_data_next[197] : sha_core_block[197];   // sha_top.v(246)
    assign n1327 = sha_state_read_data ? sha_core_block_read_data_next[196] : sha_core_block[196];   // sha_top.v(246)
    assign n1328 = sha_state_read_data ? sha_core_block_read_data_next[195] : sha_core_block[195];   // sha_top.v(246)
    assign n1329 = sha_state_read_data ? sha_core_block_read_data_next[194] : sha_core_block[194];   // sha_top.v(246)
    assign n1330 = sha_state_read_data ? sha_core_block_read_data_next[193] : sha_core_block[193];   // sha_top.v(246)
    assign n1331 = sha_state_read_data ? sha_core_block_read_data_next[192] : sha_core_block[192];   // sha_top.v(246)
    assign n1332 = sha_state_read_data ? sha_core_block_read_data_next[191] : sha_core_block[191];   // sha_top.v(246)
    assign n1333 = sha_state_read_data ? sha_core_block_read_data_next[190] : sha_core_block[190];   // sha_top.v(246)
    assign n1334 = sha_state_read_data ? sha_core_block_read_data_next[189] : sha_core_block[189];   // sha_top.v(246)
    assign n1335 = sha_state_read_data ? sha_core_block_read_data_next[188] : sha_core_block[188];   // sha_top.v(246)
    assign n1336 = sha_state_read_data ? sha_core_block_read_data_next[187] : sha_core_block[187];   // sha_top.v(246)
    assign n1337 = sha_state_read_data ? sha_core_block_read_data_next[186] : sha_core_block[186];   // sha_top.v(246)
    assign n1338 = sha_state_read_data ? sha_core_block_read_data_next[185] : sha_core_block[185];   // sha_top.v(246)
    assign n1339 = sha_state_read_data ? sha_core_block_read_data_next[184] : sha_core_block[184];   // sha_top.v(246)
    assign n1340 = sha_state_read_data ? sha_core_block_read_data_next[183] : sha_core_block[183];   // sha_top.v(246)
    assign n1341 = sha_state_read_data ? sha_core_block_read_data_next[182] : sha_core_block[182];   // sha_top.v(246)
    assign n1342 = sha_state_read_data ? sha_core_block_read_data_next[181] : sha_core_block[181];   // sha_top.v(246)
    assign n1343 = sha_state_read_data ? sha_core_block_read_data_next[180] : sha_core_block[180];   // sha_top.v(246)
    assign n1344 = sha_state_read_data ? sha_core_block_read_data_next[179] : sha_core_block[179];   // sha_top.v(246)
    assign n1345 = sha_state_read_data ? sha_core_block_read_data_next[178] : sha_core_block[178];   // sha_top.v(246)
    assign n1346 = sha_state_read_data ? sha_core_block_read_data_next[177] : sha_core_block[177];   // sha_top.v(246)
    assign n1347 = sha_state_read_data ? sha_core_block_read_data_next[176] : sha_core_block[176];   // sha_top.v(246)
    assign n1348 = sha_state_read_data ? sha_core_block_read_data_next[175] : sha_core_block[175];   // sha_top.v(246)
    assign n1349 = sha_state_read_data ? sha_core_block_read_data_next[174] : sha_core_block[174];   // sha_top.v(246)
    assign n1350 = sha_state_read_data ? sha_core_block_read_data_next[173] : sha_core_block[173];   // sha_top.v(246)
    assign n1351 = sha_state_read_data ? sha_core_block_read_data_next[172] : sha_core_block[172];   // sha_top.v(246)
    assign n1352 = sha_state_read_data ? sha_core_block_read_data_next[171] : sha_core_block[171];   // sha_top.v(246)
    assign n1353 = sha_state_read_data ? sha_core_block_read_data_next[170] : sha_core_block[170];   // sha_top.v(246)
    assign n1354 = sha_state_read_data ? sha_core_block_read_data_next[169] : sha_core_block[169];   // sha_top.v(246)
    assign n1355 = sha_state_read_data ? sha_core_block_read_data_next[168] : sha_core_block[168];   // sha_top.v(246)
    assign n1356 = sha_state_read_data ? sha_core_block_read_data_next[167] : sha_core_block[167];   // sha_top.v(246)
    assign n1357 = sha_state_read_data ? sha_core_block_read_data_next[166] : sha_core_block[166];   // sha_top.v(246)
    assign n1358 = sha_state_read_data ? sha_core_block_read_data_next[165] : sha_core_block[165];   // sha_top.v(246)
    assign n1359 = sha_state_read_data ? sha_core_block_read_data_next[164] : sha_core_block[164];   // sha_top.v(246)
    assign n1360 = sha_state_read_data ? sha_core_block_read_data_next[163] : sha_core_block[163];   // sha_top.v(246)
    assign n1361 = sha_state_read_data ? sha_core_block_read_data_next[162] : sha_core_block[162];   // sha_top.v(246)
    assign n1362 = sha_state_read_data ? sha_core_block_read_data_next[161] : sha_core_block[161];   // sha_top.v(246)
    assign n1363 = sha_state_read_data ? sha_core_block_read_data_next[160] : sha_core_block[160];   // sha_top.v(246)
    assign n1364 = sha_state_read_data ? sha_core_block_read_data_next[159] : sha_core_block[159];   // sha_top.v(246)
    assign n1365 = sha_state_read_data ? sha_core_block_read_data_next[158] : sha_core_block[158];   // sha_top.v(246)
    assign n1366 = sha_state_read_data ? sha_core_block_read_data_next[157] : sha_core_block[157];   // sha_top.v(246)
    assign n1367 = sha_state_read_data ? sha_core_block_read_data_next[156] : sha_core_block[156];   // sha_top.v(246)
    assign n1368 = sha_state_read_data ? sha_core_block_read_data_next[155] : sha_core_block[155];   // sha_top.v(246)
    assign n1369 = sha_state_read_data ? sha_core_block_read_data_next[154] : sha_core_block[154];   // sha_top.v(246)
    assign n1370 = sha_state_read_data ? sha_core_block_read_data_next[153] : sha_core_block[153];   // sha_top.v(246)
    assign n1371 = sha_state_read_data ? sha_core_block_read_data_next[152] : sha_core_block[152];   // sha_top.v(246)
    assign n1372 = sha_state_read_data ? sha_core_block_read_data_next[151] : sha_core_block[151];   // sha_top.v(246)
    assign n1373 = sha_state_read_data ? sha_core_block_read_data_next[150] : sha_core_block[150];   // sha_top.v(246)
    assign n1374 = sha_state_read_data ? sha_core_block_read_data_next[149] : sha_core_block[149];   // sha_top.v(246)
    assign n1375 = sha_state_read_data ? sha_core_block_read_data_next[148] : sha_core_block[148];   // sha_top.v(246)
    assign n1376 = sha_state_read_data ? sha_core_block_read_data_next[147] : sha_core_block[147];   // sha_top.v(246)
    assign n1377 = sha_state_read_data ? sha_core_block_read_data_next[146] : sha_core_block[146];   // sha_top.v(246)
    assign n1378 = sha_state_read_data ? sha_core_block_read_data_next[145] : sha_core_block[145];   // sha_top.v(246)
    assign n1379 = sha_state_read_data ? sha_core_block_read_data_next[144] : sha_core_block[144];   // sha_top.v(246)
    assign n1380 = sha_state_read_data ? sha_core_block_read_data_next[143] : sha_core_block[143];   // sha_top.v(246)
    assign n1381 = sha_state_read_data ? sha_core_block_read_data_next[142] : sha_core_block[142];   // sha_top.v(246)
    assign n1382 = sha_state_read_data ? sha_core_block_read_data_next[141] : sha_core_block[141];   // sha_top.v(246)
    assign n1383 = sha_state_read_data ? sha_core_block_read_data_next[140] : sha_core_block[140];   // sha_top.v(246)
    assign n1384 = sha_state_read_data ? sha_core_block_read_data_next[139] : sha_core_block[139];   // sha_top.v(246)
    assign n1385 = sha_state_read_data ? sha_core_block_read_data_next[138] : sha_core_block[138];   // sha_top.v(246)
    assign n1386 = sha_state_read_data ? sha_core_block_read_data_next[137] : sha_core_block[137];   // sha_top.v(246)
    assign n1387 = sha_state_read_data ? sha_core_block_read_data_next[136] : sha_core_block[136];   // sha_top.v(246)
    assign n1388 = sha_state_read_data ? sha_core_block_read_data_next[135] : sha_core_block[135];   // sha_top.v(246)
    assign n1389 = sha_state_read_data ? sha_core_block_read_data_next[134] : sha_core_block[134];   // sha_top.v(246)
    assign n1390 = sha_state_read_data ? sha_core_block_read_data_next[133] : sha_core_block[133];   // sha_top.v(246)
    assign n1391 = sha_state_read_data ? sha_core_block_read_data_next[132] : sha_core_block[132];   // sha_top.v(246)
    assign n1392 = sha_state_read_data ? sha_core_block_read_data_next[131] : sha_core_block[131];   // sha_top.v(246)
    assign n1393 = sha_state_read_data ? sha_core_block_read_data_next[130] : sha_core_block[130];   // sha_top.v(246)
    assign n1394 = sha_state_read_data ? sha_core_block_read_data_next[129] : sha_core_block[129];   // sha_top.v(246)
    assign n1395 = sha_state_read_data ? sha_core_block_read_data_next[128] : sha_core_block[128];   // sha_top.v(246)
    assign n1396 = sha_state_read_data ? sha_core_block_read_data_next[127] : sha_core_block[127];   // sha_top.v(246)
    assign n1397 = sha_state_read_data ? sha_core_block_read_data_next[126] : sha_core_block[126];   // sha_top.v(246)
    assign n1398 = sha_state_read_data ? sha_core_block_read_data_next[125] : sha_core_block[125];   // sha_top.v(246)
    assign n1399 = sha_state_read_data ? sha_core_block_read_data_next[124] : sha_core_block[124];   // sha_top.v(246)
    assign n1400 = sha_state_read_data ? sha_core_block_read_data_next[123] : sha_core_block[123];   // sha_top.v(246)
    assign n1401 = sha_state_read_data ? sha_core_block_read_data_next[122] : sha_core_block[122];   // sha_top.v(246)
    assign n1402 = sha_state_read_data ? sha_core_block_read_data_next[121] : sha_core_block[121];   // sha_top.v(246)
    assign n1403 = sha_state_read_data ? sha_core_block_read_data_next[120] : sha_core_block[120];   // sha_top.v(246)
    assign n1404 = sha_state_read_data ? sha_core_block_read_data_next[119] : sha_core_block[119];   // sha_top.v(246)
    assign n1405 = sha_state_read_data ? sha_core_block_read_data_next[118] : sha_core_block[118];   // sha_top.v(246)
    assign n1406 = sha_state_read_data ? sha_core_block_read_data_next[117] : sha_core_block[117];   // sha_top.v(246)
    assign n1407 = sha_state_read_data ? sha_core_block_read_data_next[116] : sha_core_block[116];   // sha_top.v(246)
    assign n1408 = sha_state_read_data ? sha_core_block_read_data_next[115] : sha_core_block[115];   // sha_top.v(246)
    assign n1409 = sha_state_read_data ? sha_core_block_read_data_next[114] : sha_core_block[114];   // sha_top.v(246)
    assign n1410 = sha_state_read_data ? sha_core_block_read_data_next[113] : sha_core_block[113];   // sha_top.v(246)
    assign n1411 = sha_state_read_data ? sha_core_block_read_data_next[112] : sha_core_block[112];   // sha_top.v(246)
    assign n1412 = sha_state_read_data ? sha_core_block_read_data_next[111] : sha_core_block[111];   // sha_top.v(246)
    assign n1413 = sha_state_read_data ? sha_core_block_read_data_next[110] : sha_core_block[110];   // sha_top.v(246)
    assign n1414 = sha_state_read_data ? sha_core_block_read_data_next[109] : sha_core_block[109];   // sha_top.v(246)
    assign n1415 = sha_state_read_data ? sha_core_block_read_data_next[108] : sha_core_block[108];   // sha_top.v(246)
    assign n1416 = sha_state_read_data ? sha_core_block_read_data_next[107] : sha_core_block[107];   // sha_top.v(246)
    assign n1417 = sha_state_read_data ? sha_core_block_read_data_next[106] : sha_core_block[106];   // sha_top.v(246)
    assign n1418 = sha_state_read_data ? sha_core_block_read_data_next[105] : sha_core_block[105];   // sha_top.v(246)
    assign n1419 = sha_state_read_data ? sha_core_block_read_data_next[104] : sha_core_block[104];   // sha_top.v(246)
    assign n1420 = sha_state_read_data ? sha_core_block_read_data_next[103] : sha_core_block[103];   // sha_top.v(246)
    assign n1421 = sha_state_read_data ? sha_core_block_read_data_next[102] : sha_core_block[102];   // sha_top.v(246)
    assign n1422 = sha_state_read_data ? sha_core_block_read_data_next[101] : sha_core_block[101];   // sha_top.v(246)
    assign n1423 = sha_state_read_data ? sha_core_block_read_data_next[100] : sha_core_block[100];   // sha_top.v(246)
    assign n1424 = sha_state_read_data ? sha_core_block_read_data_next[99] : sha_core_block[99];   // sha_top.v(246)
    assign n1425 = sha_state_read_data ? sha_core_block_read_data_next[98] : sha_core_block[98];   // sha_top.v(246)
    assign n1426 = sha_state_read_data ? sha_core_block_read_data_next[97] : sha_core_block[97];   // sha_top.v(246)
    assign n1427 = sha_state_read_data ? sha_core_block_read_data_next[96] : sha_core_block[96];   // sha_top.v(246)
    assign n1428 = sha_state_read_data ? sha_core_block_read_data_next[95] : sha_core_block[95];   // sha_top.v(246)
    assign n1429 = sha_state_read_data ? sha_core_block_read_data_next[94] : sha_core_block[94];   // sha_top.v(246)
    assign n1430 = sha_state_read_data ? sha_core_block_read_data_next[93] : sha_core_block[93];   // sha_top.v(246)
    assign n1431 = sha_state_read_data ? sha_core_block_read_data_next[92] : sha_core_block[92];   // sha_top.v(246)
    assign n1432 = sha_state_read_data ? sha_core_block_read_data_next[91] : sha_core_block[91];   // sha_top.v(246)
    assign n1433 = sha_state_read_data ? sha_core_block_read_data_next[90] : sha_core_block[90];   // sha_top.v(246)
    assign n1434 = sha_state_read_data ? sha_core_block_read_data_next[89] : sha_core_block[89];   // sha_top.v(246)
    assign n1435 = sha_state_read_data ? sha_core_block_read_data_next[88] : sha_core_block[88];   // sha_top.v(246)
    assign n1436 = sha_state_read_data ? sha_core_block_read_data_next[87] : sha_core_block[87];   // sha_top.v(246)
    assign n1437 = sha_state_read_data ? sha_core_block_read_data_next[86] : sha_core_block[86];   // sha_top.v(246)
    assign n1438 = sha_state_read_data ? sha_core_block_read_data_next[85] : sha_core_block[85];   // sha_top.v(246)
    assign n1439 = sha_state_read_data ? sha_core_block_read_data_next[84] : sha_core_block[84];   // sha_top.v(246)
    assign n1440 = sha_state_read_data ? sha_core_block_read_data_next[83] : sha_core_block[83];   // sha_top.v(246)
    assign n1441 = sha_state_read_data ? sha_core_block_read_data_next[82] : sha_core_block[82];   // sha_top.v(246)
    assign n1442 = sha_state_read_data ? sha_core_block_read_data_next[81] : sha_core_block[81];   // sha_top.v(246)
    assign n1443 = sha_state_read_data ? sha_core_block_read_data_next[80] : sha_core_block[80];   // sha_top.v(246)
    assign n1444 = sha_state_read_data ? sha_core_block_read_data_next[79] : sha_core_block[79];   // sha_top.v(246)
    assign n1445 = sha_state_read_data ? sha_core_block_read_data_next[78] : sha_core_block[78];   // sha_top.v(246)
    assign n1446 = sha_state_read_data ? sha_core_block_read_data_next[77] : sha_core_block[77];   // sha_top.v(246)
    assign n1447 = sha_state_read_data ? sha_core_block_read_data_next[76] : sha_core_block[76];   // sha_top.v(246)
    assign n1448 = sha_state_read_data ? sha_core_block_read_data_next[75] : sha_core_block[75];   // sha_top.v(246)
    assign n1449 = sha_state_read_data ? sha_core_block_read_data_next[74] : sha_core_block[74];   // sha_top.v(246)
    assign n1450 = sha_state_read_data ? sha_core_block_read_data_next[73] : sha_core_block[73];   // sha_top.v(246)
    assign n1451 = sha_state_read_data ? sha_core_block_read_data_next[72] : sha_core_block[72];   // sha_top.v(246)
    assign n1452 = sha_state_read_data ? sha_core_block_read_data_next[71] : sha_core_block[71];   // sha_top.v(246)
    assign n1453 = sha_state_read_data ? sha_core_block_read_data_next[70] : sha_core_block[70];   // sha_top.v(246)
    assign n1454 = sha_state_read_data ? sha_core_block_read_data_next[69] : sha_core_block[69];   // sha_top.v(246)
    assign n1455 = sha_state_read_data ? sha_core_block_read_data_next[68] : sha_core_block[68];   // sha_top.v(246)
    assign n1456 = sha_state_read_data ? sha_core_block_read_data_next[67] : sha_core_block[67];   // sha_top.v(246)
    assign n1457 = sha_state_read_data ? sha_core_block_read_data_next[66] : sha_core_block[66];   // sha_top.v(246)
    assign n1458 = sha_state_read_data ? sha_core_block_read_data_next[65] : sha_core_block[65];   // sha_top.v(246)
    assign n1459 = sha_state_read_data ? sha_core_block_read_data_next[64] : sha_core_block[64];   // sha_top.v(246)
    assign n1460 = sha_state_read_data ? sha_core_block_read_data_next[63] : sha_core_block[63];   // sha_top.v(246)
    assign n1461 = sha_state_read_data ? sha_core_block_read_data_next[62] : sha_core_block[62];   // sha_top.v(246)
    assign n1462 = sha_state_read_data ? sha_core_block_read_data_next[61] : sha_core_block[61];   // sha_top.v(246)
    assign n1463 = sha_state_read_data ? sha_core_block_read_data_next[60] : sha_core_block[60];   // sha_top.v(246)
    assign n1464 = sha_state_read_data ? sha_core_block_read_data_next[59] : sha_core_block[59];   // sha_top.v(246)
    assign n1465 = sha_state_read_data ? sha_core_block_read_data_next[58] : sha_core_block[58];   // sha_top.v(246)
    assign n1466 = sha_state_read_data ? sha_core_block_read_data_next[57] : sha_core_block[57];   // sha_top.v(246)
    assign n1467 = sha_state_read_data ? sha_core_block_read_data_next[56] : sha_core_block[56];   // sha_top.v(246)
    assign n1468 = sha_state_read_data ? sha_core_block_read_data_next[55] : sha_core_block[55];   // sha_top.v(246)
    assign n1469 = sha_state_read_data ? sha_core_block_read_data_next[54] : sha_core_block[54];   // sha_top.v(246)
    assign n1470 = sha_state_read_data ? sha_core_block_read_data_next[53] : sha_core_block[53];   // sha_top.v(246)
    assign n1471 = sha_state_read_data ? sha_core_block_read_data_next[52] : sha_core_block[52];   // sha_top.v(246)
    assign n1472 = sha_state_read_data ? sha_core_block_read_data_next[51] : sha_core_block[51];   // sha_top.v(246)
    assign n1473 = sha_state_read_data ? sha_core_block_read_data_next[50] : sha_core_block[50];   // sha_top.v(246)
    assign n1474 = sha_state_read_data ? sha_core_block_read_data_next[49] : sha_core_block[49];   // sha_top.v(246)
    assign n1475 = sha_state_read_data ? sha_core_block_read_data_next[48] : sha_core_block[48];   // sha_top.v(246)
    assign n1476 = sha_state_read_data ? sha_core_block_read_data_next[47] : sha_core_block[47];   // sha_top.v(246)
    assign n1477 = sha_state_read_data ? sha_core_block_read_data_next[46] : sha_core_block[46];   // sha_top.v(246)
    assign n1478 = sha_state_read_data ? sha_core_block_read_data_next[45] : sha_core_block[45];   // sha_top.v(246)
    assign n1479 = sha_state_read_data ? sha_core_block_read_data_next[44] : sha_core_block[44];   // sha_top.v(246)
    assign n1480 = sha_state_read_data ? sha_core_block_read_data_next[43] : sha_core_block[43];   // sha_top.v(246)
    assign n1481 = sha_state_read_data ? sha_core_block_read_data_next[42] : sha_core_block[42];   // sha_top.v(246)
    assign n1482 = sha_state_read_data ? sha_core_block_read_data_next[41] : sha_core_block[41];   // sha_top.v(246)
    assign n1483 = sha_state_read_data ? sha_core_block_read_data_next[40] : sha_core_block[40];   // sha_top.v(246)
    assign n1484 = sha_state_read_data ? sha_core_block_read_data_next[39] : sha_core_block[39];   // sha_top.v(246)
    assign n1485 = sha_state_read_data ? sha_core_block_read_data_next[38] : sha_core_block[38];   // sha_top.v(246)
    assign n1486 = sha_state_read_data ? sha_core_block_read_data_next[37] : sha_core_block[37];   // sha_top.v(246)
    assign n1487 = sha_state_read_data ? sha_core_block_read_data_next[36] : sha_core_block[36];   // sha_top.v(246)
    assign n1488 = sha_state_read_data ? sha_core_block_read_data_next[35] : sha_core_block[35];   // sha_top.v(246)
    assign n1489 = sha_state_read_data ? sha_core_block_read_data_next[34] : sha_core_block[34];   // sha_top.v(246)
    assign n1490 = sha_state_read_data ? sha_core_block_read_data_next[33] : sha_core_block[33];   // sha_top.v(246)
    assign n1491 = sha_state_read_data ? sha_core_block_read_data_next[32] : sha_core_block[32];   // sha_top.v(246)
    assign n1492 = sha_state_read_data ? sha_core_block_read_data_next[31] : sha_core_block[31];   // sha_top.v(246)
    assign n1493 = sha_state_read_data ? sha_core_block_read_data_next[30] : sha_core_block[30];   // sha_top.v(246)
    assign n1494 = sha_state_read_data ? sha_core_block_read_data_next[29] : sha_core_block[29];   // sha_top.v(246)
    assign n1495 = sha_state_read_data ? sha_core_block_read_data_next[28] : sha_core_block[28];   // sha_top.v(246)
    assign n1496 = sha_state_read_data ? sha_core_block_read_data_next[27] : sha_core_block[27];   // sha_top.v(246)
    assign n1497 = sha_state_read_data ? sha_core_block_read_data_next[26] : sha_core_block[26];   // sha_top.v(246)
    assign n1498 = sha_state_read_data ? sha_core_block_read_data_next[25] : sha_core_block[25];   // sha_top.v(246)
    assign n1499 = sha_state_read_data ? sha_core_block_read_data_next[24] : sha_core_block[24];   // sha_top.v(246)
    assign n1500 = sha_state_read_data ? sha_core_block_read_data_next[23] : sha_core_block[23];   // sha_top.v(246)
    assign n1501 = sha_state_read_data ? sha_core_block_read_data_next[22] : sha_core_block[22];   // sha_top.v(246)
    assign n1502 = sha_state_read_data ? sha_core_block_read_data_next[21] : sha_core_block[21];   // sha_top.v(246)
    assign n1503 = sha_state_read_data ? sha_core_block_read_data_next[20] : sha_core_block[20];   // sha_top.v(246)
    assign n1504 = sha_state_read_data ? sha_core_block_read_data_next[19] : sha_core_block[19];   // sha_top.v(246)
    assign n1505 = sha_state_read_data ? sha_core_block_read_data_next[18] : sha_core_block[18];   // sha_top.v(246)
    assign n1506 = sha_state_read_data ? sha_core_block_read_data_next[17] : sha_core_block[17];   // sha_top.v(246)
    assign n1507 = sha_state_read_data ? sha_core_block_read_data_next[16] : sha_core_block[16];   // sha_top.v(246)
    assign n1508 = sha_state_read_data ? sha_core_block_read_data_next[15] : sha_core_block[15];   // sha_top.v(246)
    assign n1509 = sha_state_read_data ? sha_core_block_read_data_next[14] : sha_core_block[14];   // sha_top.v(246)
    assign n1510 = sha_state_read_data ? sha_core_block_read_data_next[13] : sha_core_block[13];   // sha_top.v(246)
    assign n1511 = sha_state_read_data ? sha_core_block_read_data_next[12] : sha_core_block[12];   // sha_top.v(246)
    assign n1512 = sha_state_read_data ? sha_core_block_read_data_next[11] : sha_core_block[11];   // sha_top.v(246)
    assign n1513 = sha_state_read_data ? sha_core_block_read_data_next[10] : sha_core_block[10];   // sha_top.v(246)
    assign n1514 = sha_state_read_data ? sha_core_block_read_data_next[9] : sha_core_block[9];   // sha_top.v(246)
    assign n1515 = sha_state_read_data ? sha_core_block_read_data_next[8] : sha_core_block[8];   // sha_top.v(246)
    assign n1516 = sha_state_read_data ? sha_core_block_read_data_next[7] : sha_core_block[7];   // sha_top.v(246)
    assign n1517 = sha_state_read_data ? sha_core_block_read_data_next[6] : sha_core_block[6];   // sha_top.v(246)
    assign n1518 = sha_state_read_data ? sha_core_block_read_data_next[5] : sha_core_block[5];   // sha_top.v(246)
    assign n1519 = sha_state_read_data ? sha_core_block_read_data_next[4] : sha_core_block[4];   // sha_top.v(246)
    assign n1520 = sha_state_read_data ? sha_core_block_read_data_next[3] : sha_core_block[3];   // sha_top.v(246)
    assign n1521 = sha_state_read_data ? sha_core_block_read_data_next[2] : sha_core_block[2];   // sha_top.v(246)
    assign n1522 = sha_state_read_data ? sha_core_block_read_data_next[1] : sha_core_block[1];   // sha_top.v(246)
    assign n1523 = sha_state_read_data ? sha_core_block_read_data_next[0] : sha_core_block[0];   // sha_top.v(246)
    assign sha_core_block_next[511] = sha_state_idle ? 1'b0 : n1012;   // sha_top.v(246)
    assign sha_core_block_next[510] = sha_state_idle ? 1'b0 : n1013;   // sha_top.v(246)
    assign sha_core_block_next[509] = sha_state_idle ? 1'b0 : n1014;   // sha_top.v(246)
    assign sha_core_block_next[508] = sha_state_idle ? 1'b0 : n1015;   // sha_top.v(246)
    assign sha_core_block_next[507] = sha_state_idle ? 1'b0 : n1016;   // sha_top.v(246)
    assign sha_core_block_next[506] = sha_state_idle ? 1'b0 : n1017;   // sha_top.v(246)
    assign sha_core_block_next[505] = sha_state_idle ? 1'b0 : n1018;   // sha_top.v(246)
    assign sha_core_block_next[504] = sha_state_idle ? 1'b0 : n1019;   // sha_top.v(246)
    assign sha_core_block_next[503] = sha_state_idle ? 1'b0 : n1020;   // sha_top.v(246)
    assign sha_core_block_next[502] = sha_state_idle ? 1'b0 : n1021;   // sha_top.v(246)
    assign sha_core_block_next[501] = sha_state_idle ? 1'b0 : n1022;   // sha_top.v(246)
    assign sha_core_block_next[500] = sha_state_idle ? 1'b0 : n1023;   // sha_top.v(246)
    assign sha_core_block_next[499] = sha_state_idle ? 1'b0 : n1024;   // sha_top.v(246)
    assign sha_core_block_next[498] = sha_state_idle ? 1'b0 : n1025;   // sha_top.v(246)
    assign sha_core_block_next[497] = sha_state_idle ? 1'b0 : n1026;   // sha_top.v(246)
    assign sha_core_block_next[496] = sha_state_idle ? 1'b0 : n1027;   // sha_top.v(246)
    assign sha_core_block_next[495] = sha_state_idle ? 1'b0 : n1028;   // sha_top.v(246)
    assign sha_core_block_next[494] = sha_state_idle ? 1'b0 : n1029;   // sha_top.v(246)
    assign sha_core_block_next[493] = sha_state_idle ? 1'b0 : n1030;   // sha_top.v(246)
    assign sha_core_block_next[492] = sha_state_idle ? 1'b0 : n1031;   // sha_top.v(246)
    assign sha_core_block_next[491] = sha_state_idle ? 1'b0 : n1032;   // sha_top.v(246)
    assign sha_core_block_next[490] = sha_state_idle ? 1'b0 : n1033;   // sha_top.v(246)
    assign sha_core_block_next[489] = sha_state_idle ? 1'b0 : n1034;   // sha_top.v(246)
    assign sha_core_block_next[488] = sha_state_idle ? 1'b0 : n1035;   // sha_top.v(246)
    assign sha_core_block_next[487] = sha_state_idle ? 1'b0 : n1036;   // sha_top.v(246)
    assign sha_core_block_next[486] = sha_state_idle ? 1'b0 : n1037;   // sha_top.v(246)
    assign sha_core_block_next[485] = sha_state_idle ? 1'b0 : n1038;   // sha_top.v(246)
    assign sha_core_block_next[484] = sha_state_idle ? 1'b0 : n1039;   // sha_top.v(246)
    assign sha_core_block_next[483] = sha_state_idle ? 1'b0 : n1040;   // sha_top.v(246)
    assign sha_core_block_next[482] = sha_state_idle ? 1'b0 : n1041;   // sha_top.v(246)
    assign sha_core_block_next[481] = sha_state_idle ? 1'b0 : n1042;   // sha_top.v(246)
    assign sha_core_block_next[480] = sha_state_idle ? 1'b0 : n1043;   // sha_top.v(246)
    assign sha_core_block_next[479] = sha_state_idle ? 1'b0 : n1044;   // sha_top.v(246)
    assign sha_core_block_next[478] = sha_state_idle ? 1'b0 : n1045;   // sha_top.v(246)
    assign sha_core_block_next[477] = sha_state_idle ? 1'b0 : n1046;   // sha_top.v(246)
    assign sha_core_block_next[476] = sha_state_idle ? 1'b0 : n1047;   // sha_top.v(246)
    assign sha_core_block_next[475] = sha_state_idle ? 1'b0 : n1048;   // sha_top.v(246)
    assign sha_core_block_next[474] = sha_state_idle ? 1'b0 : n1049;   // sha_top.v(246)
    assign sha_core_block_next[473] = sha_state_idle ? 1'b0 : n1050;   // sha_top.v(246)
    assign sha_core_block_next[472] = sha_state_idle ? 1'b0 : n1051;   // sha_top.v(246)
    assign sha_core_block_next[471] = sha_state_idle ? 1'b0 : n1052;   // sha_top.v(246)
    assign sha_core_block_next[470] = sha_state_idle ? 1'b0 : n1053;   // sha_top.v(246)
    assign sha_core_block_next[469] = sha_state_idle ? 1'b0 : n1054;   // sha_top.v(246)
    assign sha_core_block_next[468] = sha_state_idle ? 1'b0 : n1055;   // sha_top.v(246)
    assign sha_core_block_next[467] = sha_state_idle ? 1'b0 : n1056;   // sha_top.v(246)
    assign sha_core_block_next[466] = sha_state_idle ? 1'b0 : n1057;   // sha_top.v(246)
    assign sha_core_block_next[465] = sha_state_idle ? 1'b0 : n1058;   // sha_top.v(246)
    assign sha_core_block_next[464] = sha_state_idle ? 1'b0 : n1059;   // sha_top.v(246)
    assign sha_core_block_next[463] = sha_state_idle ? 1'b0 : n1060;   // sha_top.v(246)
    assign sha_core_block_next[462] = sha_state_idle ? 1'b0 : n1061;   // sha_top.v(246)
    assign sha_core_block_next[461] = sha_state_idle ? 1'b0 : n1062;   // sha_top.v(246)
    assign sha_core_block_next[460] = sha_state_idle ? 1'b0 : n1063;   // sha_top.v(246)
    assign sha_core_block_next[459] = sha_state_idle ? 1'b0 : n1064;   // sha_top.v(246)
    assign sha_core_block_next[458] = sha_state_idle ? 1'b0 : n1065;   // sha_top.v(246)
    assign sha_core_block_next[457] = sha_state_idle ? 1'b0 : n1066;   // sha_top.v(246)
    assign sha_core_block_next[456] = sha_state_idle ? 1'b0 : n1067;   // sha_top.v(246)
    assign sha_core_block_next[455] = sha_state_idle ? 1'b0 : n1068;   // sha_top.v(246)
    assign sha_core_block_next[454] = sha_state_idle ? 1'b0 : n1069;   // sha_top.v(246)
    assign sha_core_block_next[453] = sha_state_idle ? 1'b0 : n1070;   // sha_top.v(246)
    assign sha_core_block_next[452] = sha_state_idle ? 1'b0 : n1071;   // sha_top.v(246)
    assign sha_core_block_next[451] = sha_state_idle ? 1'b0 : n1072;   // sha_top.v(246)
    assign sha_core_block_next[450] = sha_state_idle ? 1'b0 : n1073;   // sha_top.v(246)
    assign sha_core_block_next[449] = sha_state_idle ? 1'b0 : n1074;   // sha_top.v(246)
    assign sha_core_block_next[448] = sha_state_idle ? 1'b0 : n1075;   // sha_top.v(246)
    assign sha_core_block_next[447] = sha_state_idle ? 1'b0 : n1076;   // sha_top.v(246)
    assign sha_core_block_next[446] = sha_state_idle ? 1'b0 : n1077;   // sha_top.v(246)
    assign sha_core_block_next[445] = sha_state_idle ? 1'b0 : n1078;   // sha_top.v(246)
    assign sha_core_block_next[444] = sha_state_idle ? 1'b0 : n1079;   // sha_top.v(246)
    assign sha_core_block_next[443] = sha_state_idle ? 1'b0 : n1080;   // sha_top.v(246)
    assign sha_core_block_next[442] = sha_state_idle ? 1'b0 : n1081;   // sha_top.v(246)
    assign sha_core_block_next[441] = sha_state_idle ? 1'b0 : n1082;   // sha_top.v(246)
    assign sha_core_block_next[440] = sha_state_idle ? 1'b0 : n1083;   // sha_top.v(246)
    assign sha_core_block_next[439] = sha_state_idle ? 1'b0 : n1084;   // sha_top.v(246)
    assign sha_core_block_next[438] = sha_state_idle ? 1'b0 : n1085;   // sha_top.v(246)
    assign sha_core_block_next[437] = sha_state_idle ? 1'b0 : n1086;   // sha_top.v(246)
    assign sha_core_block_next[436] = sha_state_idle ? 1'b0 : n1087;   // sha_top.v(246)
    assign sha_core_block_next[435] = sha_state_idle ? 1'b0 : n1088;   // sha_top.v(246)
    assign sha_core_block_next[434] = sha_state_idle ? 1'b0 : n1089;   // sha_top.v(246)
    assign sha_core_block_next[433] = sha_state_idle ? 1'b0 : n1090;   // sha_top.v(246)
    assign sha_core_block_next[432] = sha_state_idle ? 1'b0 : n1091;   // sha_top.v(246)
    assign sha_core_block_next[431] = sha_state_idle ? 1'b0 : n1092;   // sha_top.v(246)
    assign sha_core_block_next[430] = sha_state_idle ? 1'b0 : n1093;   // sha_top.v(246)
    assign sha_core_block_next[429] = sha_state_idle ? 1'b0 : n1094;   // sha_top.v(246)
    assign sha_core_block_next[428] = sha_state_idle ? 1'b0 : n1095;   // sha_top.v(246)
    assign sha_core_block_next[427] = sha_state_idle ? 1'b0 : n1096;   // sha_top.v(246)
    assign sha_core_block_next[426] = sha_state_idle ? 1'b0 : n1097;   // sha_top.v(246)
    assign sha_core_block_next[425] = sha_state_idle ? 1'b0 : n1098;   // sha_top.v(246)
    assign sha_core_block_next[424] = sha_state_idle ? 1'b0 : n1099;   // sha_top.v(246)
    assign sha_core_block_next[423] = sha_state_idle ? 1'b0 : n1100;   // sha_top.v(246)
    assign sha_core_block_next[422] = sha_state_idle ? 1'b0 : n1101;   // sha_top.v(246)
    assign sha_core_block_next[421] = sha_state_idle ? 1'b0 : n1102;   // sha_top.v(246)
    assign sha_core_block_next[420] = sha_state_idle ? 1'b0 : n1103;   // sha_top.v(246)
    assign sha_core_block_next[419] = sha_state_idle ? 1'b0 : n1104;   // sha_top.v(246)
    assign sha_core_block_next[418] = sha_state_idle ? 1'b0 : n1105;   // sha_top.v(246)
    assign sha_core_block_next[417] = sha_state_idle ? 1'b0 : n1106;   // sha_top.v(246)
    assign sha_core_block_next[416] = sha_state_idle ? 1'b0 : n1107;   // sha_top.v(246)
    assign sha_core_block_next[415] = sha_state_idle ? 1'b0 : n1108;   // sha_top.v(246)
    assign sha_core_block_next[414] = sha_state_idle ? 1'b0 : n1109;   // sha_top.v(246)
    assign sha_core_block_next[413] = sha_state_idle ? 1'b0 : n1110;   // sha_top.v(246)
    assign sha_core_block_next[412] = sha_state_idle ? 1'b0 : n1111;   // sha_top.v(246)
    assign sha_core_block_next[411] = sha_state_idle ? 1'b0 : n1112;   // sha_top.v(246)
    assign sha_core_block_next[410] = sha_state_idle ? 1'b0 : n1113;   // sha_top.v(246)
    assign sha_core_block_next[409] = sha_state_idle ? 1'b0 : n1114;   // sha_top.v(246)
    assign sha_core_block_next[408] = sha_state_idle ? 1'b0 : n1115;   // sha_top.v(246)
    assign sha_core_block_next[407] = sha_state_idle ? 1'b0 : n1116;   // sha_top.v(246)
    assign sha_core_block_next[406] = sha_state_idle ? 1'b0 : n1117;   // sha_top.v(246)
    assign sha_core_block_next[405] = sha_state_idle ? 1'b0 : n1118;   // sha_top.v(246)
    assign sha_core_block_next[404] = sha_state_idle ? 1'b0 : n1119;   // sha_top.v(246)
    assign sha_core_block_next[403] = sha_state_idle ? 1'b0 : n1120;   // sha_top.v(246)
    assign sha_core_block_next[402] = sha_state_idle ? 1'b0 : n1121;   // sha_top.v(246)
    assign sha_core_block_next[401] = sha_state_idle ? 1'b0 : n1122;   // sha_top.v(246)
    assign sha_core_block_next[400] = sha_state_idle ? 1'b0 : n1123;   // sha_top.v(246)
    assign sha_core_block_next[399] = sha_state_idle ? 1'b0 : n1124;   // sha_top.v(246)
    assign sha_core_block_next[398] = sha_state_idle ? 1'b0 : n1125;   // sha_top.v(246)
    assign sha_core_block_next[397] = sha_state_idle ? 1'b0 : n1126;   // sha_top.v(246)
    assign sha_core_block_next[396] = sha_state_idle ? 1'b0 : n1127;   // sha_top.v(246)
    assign sha_core_block_next[395] = sha_state_idle ? 1'b0 : n1128;   // sha_top.v(246)
    assign sha_core_block_next[394] = sha_state_idle ? 1'b0 : n1129;   // sha_top.v(246)
    assign sha_core_block_next[393] = sha_state_idle ? 1'b0 : n1130;   // sha_top.v(246)
    assign sha_core_block_next[392] = sha_state_idle ? 1'b0 : n1131;   // sha_top.v(246)
    assign sha_core_block_next[391] = sha_state_idle ? 1'b0 : n1132;   // sha_top.v(246)
    assign sha_core_block_next[390] = sha_state_idle ? 1'b0 : n1133;   // sha_top.v(246)
    assign sha_core_block_next[389] = sha_state_idle ? 1'b0 : n1134;   // sha_top.v(246)
    assign sha_core_block_next[388] = sha_state_idle ? 1'b0 : n1135;   // sha_top.v(246)
    assign sha_core_block_next[387] = sha_state_idle ? 1'b0 : n1136;   // sha_top.v(246)
    assign sha_core_block_next[386] = sha_state_idle ? 1'b0 : n1137;   // sha_top.v(246)
    assign sha_core_block_next[385] = sha_state_idle ? 1'b0 : n1138;   // sha_top.v(246)
    assign sha_core_block_next[384] = sha_state_idle ? 1'b0 : n1139;   // sha_top.v(246)
    assign sha_core_block_next[383] = sha_state_idle ? 1'b0 : n1140;   // sha_top.v(246)
    assign sha_core_block_next[382] = sha_state_idle ? 1'b0 : n1141;   // sha_top.v(246)
    assign sha_core_block_next[381] = sha_state_idle ? 1'b0 : n1142;   // sha_top.v(246)
    assign sha_core_block_next[380] = sha_state_idle ? 1'b0 : n1143;   // sha_top.v(246)
    assign sha_core_block_next[379] = sha_state_idle ? 1'b0 : n1144;   // sha_top.v(246)
    assign sha_core_block_next[378] = sha_state_idle ? 1'b0 : n1145;   // sha_top.v(246)
    assign sha_core_block_next[377] = sha_state_idle ? 1'b0 : n1146;   // sha_top.v(246)
    assign sha_core_block_next[376] = sha_state_idle ? 1'b0 : n1147;   // sha_top.v(246)
    assign sha_core_block_next[375] = sha_state_idle ? 1'b0 : n1148;   // sha_top.v(246)
    assign sha_core_block_next[374] = sha_state_idle ? 1'b0 : n1149;   // sha_top.v(246)
    assign sha_core_block_next[373] = sha_state_idle ? 1'b0 : n1150;   // sha_top.v(246)
    assign sha_core_block_next[372] = sha_state_idle ? 1'b0 : n1151;   // sha_top.v(246)
    assign sha_core_block_next[371] = sha_state_idle ? 1'b0 : n1152;   // sha_top.v(246)
    assign sha_core_block_next[370] = sha_state_idle ? 1'b0 : n1153;   // sha_top.v(246)
    assign sha_core_block_next[369] = sha_state_idle ? 1'b0 : n1154;   // sha_top.v(246)
    assign sha_core_block_next[368] = sha_state_idle ? 1'b0 : n1155;   // sha_top.v(246)
    assign sha_core_block_next[367] = sha_state_idle ? 1'b0 : n1156;   // sha_top.v(246)
    assign sha_core_block_next[366] = sha_state_idle ? 1'b0 : n1157;   // sha_top.v(246)
    assign sha_core_block_next[365] = sha_state_idle ? 1'b0 : n1158;   // sha_top.v(246)
    assign sha_core_block_next[364] = sha_state_idle ? 1'b0 : n1159;   // sha_top.v(246)
    assign sha_core_block_next[363] = sha_state_idle ? 1'b0 : n1160;   // sha_top.v(246)
    assign sha_core_block_next[362] = sha_state_idle ? 1'b0 : n1161;   // sha_top.v(246)
    assign sha_core_block_next[361] = sha_state_idle ? 1'b0 : n1162;   // sha_top.v(246)
    assign sha_core_block_next[360] = sha_state_idle ? 1'b0 : n1163;   // sha_top.v(246)
    assign sha_core_block_next[359] = sha_state_idle ? 1'b0 : n1164;   // sha_top.v(246)
    assign sha_core_block_next[358] = sha_state_idle ? 1'b0 : n1165;   // sha_top.v(246)
    assign sha_core_block_next[357] = sha_state_idle ? 1'b0 : n1166;   // sha_top.v(246)
    assign sha_core_block_next[356] = sha_state_idle ? 1'b0 : n1167;   // sha_top.v(246)
    assign sha_core_block_next[355] = sha_state_idle ? 1'b0 : n1168;   // sha_top.v(246)
    assign sha_core_block_next[354] = sha_state_idle ? 1'b0 : n1169;   // sha_top.v(246)
    assign sha_core_block_next[353] = sha_state_idle ? 1'b0 : n1170;   // sha_top.v(246)
    assign sha_core_block_next[352] = sha_state_idle ? 1'b0 : n1171;   // sha_top.v(246)
    assign sha_core_block_next[351] = sha_state_idle ? 1'b0 : n1172;   // sha_top.v(246)
    assign sha_core_block_next[350] = sha_state_idle ? 1'b0 : n1173;   // sha_top.v(246)
    assign sha_core_block_next[349] = sha_state_idle ? 1'b0 : n1174;   // sha_top.v(246)
    assign sha_core_block_next[348] = sha_state_idle ? 1'b0 : n1175;   // sha_top.v(246)
    assign sha_core_block_next[347] = sha_state_idle ? 1'b0 : n1176;   // sha_top.v(246)
    assign sha_core_block_next[346] = sha_state_idle ? 1'b0 : n1177;   // sha_top.v(246)
    assign sha_core_block_next[345] = sha_state_idle ? 1'b0 : n1178;   // sha_top.v(246)
    assign sha_core_block_next[344] = sha_state_idle ? 1'b0 : n1179;   // sha_top.v(246)
    assign sha_core_block_next[343] = sha_state_idle ? 1'b0 : n1180;   // sha_top.v(246)
    assign sha_core_block_next[342] = sha_state_idle ? 1'b0 : n1181;   // sha_top.v(246)
    assign sha_core_block_next[341] = sha_state_idle ? 1'b0 : n1182;   // sha_top.v(246)
    assign sha_core_block_next[340] = sha_state_idle ? 1'b0 : n1183;   // sha_top.v(246)
    assign sha_core_block_next[339] = sha_state_idle ? 1'b0 : n1184;   // sha_top.v(246)
    assign sha_core_block_next[338] = sha_state_idle ? 1'b0 : n1185;   // sha_top.v(246)
    assign sha_core_block_next[337] = sha_state_idle ? 1'b0 : n1186;   // sha_top.v(246)
    assign sha_core_block_next[336] = sha_state_idle ? 1'b0 : n1187;   // sha_top.v(246)
    assign sha_core_block_next[335] = sha_state_idle ? 1'b0 : n1188;   // sha_top.v(246)
    assign sha_core_block_next[334] = sha_state_idle ? 1'b0 : n1189;   // sha_top.v(246)
    assign sha_core_block_next[333] = sha_state_idle ? 1'b0 : n1190;   // sha_top.v(246)
    assign sha_core_block_next[332] = sha_state_idle ? 1'b0 : n1191;   // sha_top.v(246)
    assign sha_core_block_next[331] = sha_state_idle ? 1'b0 : n1192;   // sha_top.v(246)
    assign sha_core_block_next[330] = sha_state_idle ? 1'b0 : n1193;   // sha_top.v(246)
    assign sha_core_block_next[329] = sha_state_idle ? 1'b0 : n1194;   // sha_top.v(246)
    assign sha_core_block_next[328] = sha_state_idle ? 1'b0 : n1195;   // sha_top.v(246)
    assign sha_core_block_next[327] = sha_state_idle ? 1'b0 : n1196;   // sha_top.v(246)
    assign sha_core_block_next[326] = sha_state_idle ? 1'b0 : n1197;   // sha_top.v(246)
    assign sha_core_block_next[325] = sha_state_idle ? 1'b0 : n1198;   // sha_top.v(246)
    assign sha_core_block_next[324] = sha_state_idle ? 1'b0 : n1199;   // sha_top.v(246)
    assign sha_core_block_next[323] = sha_state_idle ? 1'b0 : n1200;   // sha_top.v(246)
    assign sha_core_block_next[322] = sha_state_idle ? 1'b0 : n1201;   // sha_top.v(246)
    assign sha_core_block_next[321] = sha_state_idle ? 1'b0 : n1202;   // sha_top.v(246)
    assign sha_core_block_next[320] = sha_state_idle ? 1'b0 : n1203;   // sha_top.v(246)
    assign sha_core_block_next[319] = sha_state_idle ? 1'b0 : n1204;   // sha_top.v(246)
    assign sha_core_block_next[318] = sha_state_idle ? 1'b0 : n1205;   // sha_top.v(246)
    assign sha_core_block_next[317] = sha_state_idle ? 1'b0 : n1206;   // sha_top.v(246)
    assign sha_core_block_next[316] = sha_state_idle ? 1'b0 : n1207;   // sha_top.v(246)
    assign sha_core_block_next[315] = sha_state_idle ? 1'b0 : n1208;   // sha_top.v(246)
    assign sha_core_block_next[314] = sha_state_idle ? 1'b0 : n1209;   // sha_top.v(246)
    assign sha_core_block_next[313] = sha_state_idle ? 1'b0 : n1210;   // sha_top.v(246)
    assign sha_core_block_next[312] = sha_state_idle ? 1'b0 : n1211;   // sha_top.v(246)
    assign sha_core_block_next[311] = sha_state_idle ? 1'b0 : n1212;   // sha_top.v(246)
    assign sha_core_block_next[310] = sha_state_idle ? 1'b0 : n1213;   // sha_top.v(246)
    assign sha_core_block_next[309] = sha_state_idle ? 1'b0 : n1214;   // sha_top.v(246)
    assign sha_core_block_next[308] = sha_state_idle ? 1'b0 : n1215;   // sha_top.v(246)
    assign sha_core_block_next[307] = sha_state_idle ? 1'b0 : n1216;   // sha_top.v(246)
    assign sha_core_block_next[306] = sha_state_idle ? 1'b0 : n1217;   // sha_top.v(246)
    assign sha_core_block_next[305] = sha_state_idle ? 1'b0 : n1218;   // sha_top.v(246)
    assign sha_core_block_next[304] = sha_state_idle ? 1'b0 : n1219;   // sha_top.v(246)
    assign sha_core_block_next[303] = sha_state_idle ? 1'b0 : n1220;   // sha_top.v(246)
    assign sha_core_block_next[302] = sha_state_idle ? 1'b0 : n1221;   // sha_top.v(246)
    assign sha_core_block_next[301] = sha_state_idle ? 1'b0 : n1222;   // sha_top.v(246)
    assign sha_core_block_next[300] = sha_state_idle ? 1'b0 : n1223;   // sha_top.v(246)
    assign sha_core_block_next[299] = sha_state_idle ? 1'b0 : n1224;   // sha_top.v(246)
    assign sha_core_block_next[298] = sha_state_idle ? 1'b0 : n1225;   // sha_top.v(246)
    assign sha_core_block_next[297] = sha_state_idle ? 1'b0 : n1226;   // sha_top.v(246)
    assign sha_core_block_next[296] = sha_state_idle ? 1'b0 : n1227;   // sha_top.v(246)
    assign sha_core_block_next[295] = sha_state_idle ? 1'b0 : n1228;   // sha_top.v(246)
    assign sha_core_block_next[294] = sha_state_idle ? 1'b0 : n1229;   // sha_top.v(246)
    assign sha_core_block_next[293] = sha_state_idle ? 1'b0 : n1230;   // sha_top.v(246)
    assign sha_core_block_next[292] = sha_state_idle ? 1'b0 : n1231;   // sha_top.v(246)
    assign sha_core_block_next[291] = sha_state_idle ? 1'b0 : n1232;   // sha_top.v(246)
    assign sha_core_block_next[290] = sha_state_idle ? 1'b0 : n1233;   // sha_top.v(246)
    assign sha_core_block_next[289] = sha_state_idle ? 1'b0 : n1234;   // sha_top.v(246)
    assign sha_core_block_next[288] = sha_state_idle ? 1'b0 : n1235;   // sha_top.v(246)
    assign sha_core_block_next[287] = sha_state_idle ? 1'b0 : n1236;   // sha_top.v(246)
    assign sha_core_block_next[286] = sha_state_idle ? 1'b0 : n1237;   // sha_top.v(246)
    assign sha_core_block_next[285] = sha_state_idle ? 1'b0 : n1238;   // sha_top.v(246)
    assign sha_core_block_next[284] = sha_state_idle ? 1'b0 : n1239;   // sha_top.v(246)
    assign sha_core_block_next[283] = sha_state_idle ? 1'b0 : n1240;   // sha_top.v(246)
    assign sha_core_block_next[282] = sha_state_idle ? 1'b0 : n1241;   // sha_top.v(246)
    assign sha_core_block_next[281] = sha_state_idle ? 1'b0 : n1242;   // sha_top.v(246)
    assign sha_core_block_next[280] = sha_state_idle ? 1'b0 : n1243;   // sha_top.v(246)
    assign sha_core_block_next[279] = sha_state_idle ? 1'b0 : n1244;   // sha_top.v(246)
    assign sha_core_block_next[278] = sha_state_idle ? 1'b0 : n1245;   // sha_top.v(246)
    assign sha_core_block_next[277] = sha_state_idle ? 1'b0 : n1246;   // sha_top.v(246)
    assign sha_core_block_next[276] = sha_state_idle ? 1'b0 : n1247;   // sha_top.v(246)
    assign sha_core_block_next[275] = sha_state_idle ? 1'b0 : n1248;   // sha_top.v(246)
    assign sha_core_block_next[274] = sha_state_idle ? 1'b0 : n1249;   // sha_top.v(246)
    assign sha_core_block_next[273] = sha_state_idle ? 1'b0 : n1250;   // sha_top.v(246)
    assign sha_core_block_next[272] = sha_state_idle ? 1'b0 : n1251;   // sha_top.v(246)
    assign sha_core_block_next[271] = sha_state_idle ? 1'b0 : n1252;   // sha_top.v(246)
    assign sha_core_block_next[270] = sha_state_idle ? 1'b0 : n1253;   // sha_top.v(246)
    assign sha_core_block_next[269] = sha_state_idle ? 1'b0 : n1254;   // sha_top.v(246)
    assign sha_core_block_next[268] = sha_state_idle ? 1'b0 : n1255;   // sha_top.v(246)
    assign sha_core_block_next[267] = sha_state_idle ? 1'b0 : n1256;   // sha_top.v(246)
    assign sha_core_block_next[266] = sha_state_idle ? 1'b0 : n1257;   // sha_top.v(246)
    assign sha_core_block_next[265] = sha_state_idle ? 1'b0 : n1258;   // sha_top.v(246)
    assign sha_core_block_next[264] = sha_state_idle ? 1'b0 : n1259;   // sha_top.v(246)
    assign sha_core_block_next[263] = sha_state_idle ? 1'b0 : n1260;   // sha_top.v(246)
    assign sha_core_block_next[262] = sha_state_idle ? 1'b0 : n1261;   // sha_top.v(246)
    assign sha_core_block_next[261] = sha_state_idle ? 1'b0 : n1262;   // sha_top.v(246)
    assign sha_core_block_next[260] = sha_state_idle ? 1'b0 : n1263;   // sha_top.v(246)
    assign sha_core_block_next[259] = sha_state_idle ? 1'b0 : n1264;   // sha_top.v(246)
    assign sha_core_block_next[258] = sha_state_idle ? 1'b0 : n1265;   // sha_top.v(246)
    assign sha_core_block_next[257] = sha_state_idle ? 1'b0 : n1266;   // sha_top.v(246)
    assign sha_core_block_next[256] = sha_state_idle ? 1'b0 : n1267;   // sha_top.v(246)
    assign sha_core_block_next[255] = sha_state_idle ? 1'b0 : n1268;   // sha_top.v(246)
    assign sha_core_block_next[254] = sha_state_idle ? 1'b0 : n1269;   // sha_top.v(246)
    assign sha_core_block_next[253] = sha_state_idle ? 1'b0 : n1270;   // sha_top.v(246)
    assign sha_core_block_next[252] = sha_state_idle ? 1'b0 : n1271;   // sha_top.v(246)
    assign sha_core_block_next[251] = sha_state_idle ? 1'b0 : n1272;   // sha_top.v(246)
    assign sha_core_block_next[250] = sha_state_idle ? 1'b0 : n1273;   // sha_top.v(246)
    assign sha_core_block_next[249] = sha_state_idle ? 1'b0 : n1274;   // sha_top.v(246)
    assign sha_core_block_next[248] = sha_state_idle ? 1'b0 : n1275;   // sha_top.v(246)
    assign sha_core_block_next[247] = sha_state_idle ? 1'b0 : n1276;   // sha_top.v(246)
    assign sha_core_block_next[246] = sha_state_idle ? 1'b0 : n1277;   // sha_top.v(246)
    assign sha_core_block_next[245] = sha_state_idle ? 1'b0 : n1278;   // sha_top.v(246)
    assign sha_core_block_next[244] = sha_state_idle ? 1'b0 : n1279;   // sha_top.v(246)
    assign sha_core_block_next[243] = sha_state_idle ? 1'b0 : n1280;   // sha_top.v(246)
    assign sha_core_block_next[242] = sha_state_idle ? 1'b0 : n1281;   // sha_top.v(246)
    assign sha_core_block_next[241] = sha_state_idle ? 1'b0 : n1282;   // sha_top.v(246)
    assign sha_core_block_next[240] = sha_state_idle ? 1'b0 : n1283;   // sha_top.v(246)
    assign sha_core_block_next[239] = sha_state_idle ? 1'b0 : n1284;   // sha_top.v(246)
    assign sha_core_block_next[238] = sha_state_idle ? 1'b0 : n1285;   // sha_top.v(246)
    assign sha_core_block_next[237] = sha_state_idle ? 1'b0 : n1286;   // sha_top.v(246)
    assign sha_core_block_next[236] = sha_state_idle ? 1'b0 : n1287;   // sha_top.v(246)
    assign sha_core_block_next[235] = sha_state_idle ? 1'b0 : n1288;   // sha_top.v(246)
    assign sha_core_block_next[234] = sha_state_idle ? 1'b0 : n1289;   // sha_top.v(246)
    assign sha_core_block_next[233] = sha_state_idle ? 1'b0 : n1290;   // sha_top.v(246)
    assign sha_core_block_next[232] = sha_state_idle ? 1'b0 : n1291;   // sha_top.v(246)
    assign sha_core_block_next[231] = sha_state_idle ? 1'b0 : n1292;   // sha_top.v(246)
    assign sha_core_block_next[230] = sha_state_idle ? 1'b0 : n1293;   // sha_top.v(246)
    assign sha_core_block_next[229] = sha_state_idle ? 1'b0 : n1294;   // sha_top.v(246)
    assign sha_core_block_next[228] = sha_state_idle ? 1'b0 : n1295;   // sha_top.v(246)
    assign sha_core_block_next[227] = sha_state_idle ? 1'b0 : n1296;   // sha_top.v(246)
    assign sha_core_block_next[226] = sha_state_idle ? 1'b0 : n1297;   // sha_top.v(246)
    assign sha_core_block_next[225] = sha_state_idle ? 1'b0 : n1298;   // sha_top.v(246)
    assign sha_core_block_next[224] = sha_state_idle ? 1'b0 : n1299;   // sha_top.v(246)
    assign sha_core_block_next[223] = sha_state_idle ? 1'b0 : n1300;   // sha_top.v(246)
    assign sha_core_block_next[222] = sha_state_idle ? 1'b0 : n1301;   // sha_top.v(246)
    assign sha_core_block_next[221] = sha_state_idle ? 1'b0 : n1302;   // sha_top.v(246)
    assign sha_core_block_next[220] = sha_state_idle ? 1'b0 : n1303;   // sha_top.v(246)
    assign sha_core_block_next[219] = sha_state_idle ? 1'b0 : n1304;   // sha_top.v(246)
    assign sha_core_block_next[218] = sha_state_idle ? 1'b0 : n1305;   // sha_top.v(246)
    assign sha_core_block_next[217] = sha_state_idle ? 1'b0 : n1306;   // sha_top.v(246)
    assign sha_core_block_next[216] = sha_state_idle ? 1'b0 : n1307;   // sha_top.v(246)
    assign sha_core_block_next[215] = sha_state_idle ? 1'b0 : n1308;   // sha_top.v(246)
    assign sha_core_block_next[214] = sha_state_idle ? 1'b0 : n1309;   // sha_top.v(246)
    assign sha_core_block_next[213] = sha_state_idle ? 1'b0 : n1310;   // sha_top.v(246)
    assign sha_core_block_next[212] = sha_state_idle ? 1'b0 : n1311;   // sha_top.v(246)
    assign sha_core_block_next[211] = sha_state_idle ? 1'b0 : n1312;   // sha_top.v(246)
    assign sha_core_block_next[210] = sha_state_idle ? 1'b0 : n1313;   // sha_top.v(246)
    assign sha_core_block_next[209] = sha_state_idle ? 1'b0 : n1314;   // sha_top.v(246)
    assign sha_core_block_next[208] = sha_state_idle ? 1'b0 : n1315;   // sha_top.v(246)
    assign sha_core_block_next[207] = sha_state_idle ? 1'b0 : n1316;   // sha_top.v(246)
    assign sha_core_block_next[206] = sha_state_idle ? 1'b0 : n1317;   // sha_top.v(246)
    assign sha_core_block_next[205] = sha_state_idle ? 1'b0 : n1318;   // sha_top.v(246)
    assign sha_core_block_next[204] = sha_state_idle ? 1'b0 : n1319;   // sha_top.v(246)
    assign sha_core_block_next[203] = sha_state_idle ? 1'b0 : n1320;   // sha_top.v(246)
    assign sha_core_block_next[202] = sha_state_idle ? 1'b0 : n1321;   // sha_top.v(246)
    assign sha_core_block_next[201] = sha_state_idle ? 1'b0 : n1322;   // sha_top.v(246)
    assign sha_core_block_next[200] = sha_state_idle ? 1'b0 : n1323;   // sha_top.v(246)
    assign sha_core_block_next[199] = sha_state_idle ? 1'b0 : n1324;   // sha_top.v(246)
    assign sha_core_block_next[198] = sha_state_idle ? 1'b0 : n1325;   // sha_top.v(246)
    assign sha_core_block_next[197] = sha_state_idle ? 1'b0 : n1326;   // sha_top.v(246)
    assign sha_core_block_next[196] = sha_state_idle ? 1'b0 : n1327;   // sha_top.v(246)
    assign sha_core_block_next[195] = sha_state_idle ? 1'b0 : n1328;   // sha_top.v(246)
    assign sha_core_block_next[194] = sha_state_idle ? 1'b0 : n1329;   // sha_top.v(246)
    assign sha_core_block_next[193] = sha_state_idle ? 1'b0 : n1330;   // sha_top.v(246)
    assign sha_core_block_next[192] = sha_state_idle ? 1'b0 : n1331;   // sha_top.v(246)
    assign sha_core_block_next[191] = sha_state_idle ? 1'b0 : n1332;   // sha_top.v(246)
    assign sha_core_block_next[190] = sha_state_idle ? 1'b0 : n1333;   // sha_top.v(246)
    assign sha_core_block_next[189] = sha_state_idle ? 1'b0 : n1334;   // sha_top.v(246)
    assign sha_core_block_next[188] = sha_state_idle ? 1'b0 : n1335;   // sha_top.v(246)
    assign sha_core_block_next[187] = sha_state_idle ? 1'b0 : n1336;   // sha_top.v(246)
    assign sha_core_block_next[186] = sha_state_idle ? 1'b0 : n1337;   // sha_top.v(246)
    assign sha_core_block_next[185] = sha_state_idle ? 1'b0 : n1338;   // sha_top.v(246)
    assign sha_core_block_next[184] = sha_state_idle ? 1'b0 : n1339;   // sha_top.v(246)
    assign sha_core_block_next[183] = sha_state_idle ? 1'b0 : n1340;   // sha_top.v(246)
    assign sha_core_block_next[182] = sha_state_idle ? 1'b0 : n1341;   // sha_top.v(246)
    assign sha_core_block_next[181] = sha_state_idle ? 1'b0 : n1342;   // sha_top.v(246)
    assign sha_core_block_next[180] = sha_state_idle ? 1'b0 : n1343;   // sha_top.v(246)
    assign sha_core_block_next[179] = sha_state_idle ? 1'b0 : n1344;   // sha_top.v(246)
    assign sha_core_block_next[178] = sha_state_idle ? 1'b0 : n1345;   // sha_top.v(246)
    assign sha_core_block_next[177] = sha_state_idle ? 1'b0 : n1346;   // sha_top.v(246)
    assign sha_core_block_next[176] = sha_state_idle ? 1'b0 : n1347;   // sha_top.v(246)
    assign sha_core_block_next[175] = sha_state_idle ? 1'b0 : n1348;   // sha_top.v(246)
    assign sha_core_block_next[174] = sha_state_idle ? 1'b0 : n1349;   // sha_top.v(246)
    assign sha_core_block_next[173] = sha_state_idle ? 1'b0 : n1350;   // sha_top.v(246)
    assign sha_core_block_next[172] = sha_state_idle ? 1'b0 : n1351;   // sha_top.v(246)
    assign sha_core_block_next[171] = sha_state_idle ? 1'b0 : n1352;   // sha_top.v(246)
    assign sha_core_block_next[170] = sha_state_idle ? 1'b0 : n1353;   // sha_top.v(246)
    assign sha_core_block_next[169] = sha_state_idle ? 1'b0 : n1354;   // sha_top.v(246)
    assign sha_core_block_next[168] = sha_state_idle ? 1'b0 : n1355;   // sha_top.v(246)
    assign sha_core_block_next[167] = sha_state_idle ? 1'b0 : n1356;   // sha_top.v(246)
    assign sha_core_block_next[166] = sha_state_idle ? 1'b0 : n1357;   // sha_top.v(246)
    assign sha_core_block_next[165] = sha_state_idle ? 1'b0 : n1358;   // sha_top.v(246)
    assign sha_core_block_next[164] = sha_state_idle ? 1'b0 : n1359;   // sha_top.v(246)
    assign sha_core_block_next[163] = sha_state_idle ? 1'b0 : n1360;   // sha_top.v(246)
    assign sha_core_block_next[162] = sha_state_idle ? 1'b0 : n1361;   // sha_top.v(246)
    assign sha_core_block_next[161] = sha_state_idle ? 1'b0 : n1362;   // sha_top.v(246)
    assign sha_core_block_next[160] = sha_state_idle ? 1'b0 : n1363;   // sha_top.v(246)
    assign sha_core_block_next[159] = sha_state_idle ? 1'b0 : n1364;   // sha_top.v(246)
    assign sha_core_block_next[158] = sha_state_idle ? 1'b0 : n1365;   // sha_top.v(246)
    assign sha_core_block_next[157] = sha_state_idle ? 1'b0 : n1366;   // sha_top.v(246)
    assign sha_core_block_next[156] = sha_state_idle ? 1'b0 : n1367;   // sha_top.v(246)
    assign sha_core_block_next[155] = sha_state_idle ? 1'b0 : n1368;   // sha_top.v(246)
    assign sha_core_block_next[154] = sha_state_idle ? 1'b0 : n1369;   // sha_top.v(246)
    assign sha_core_block_next[153] = sha_state_idle ? 1'b0 : n1370;   // sha_top.v(246)
    assign sha_core_block_next[152] = sha_state_idle ? 1'b0 : n1371;   // sha_top.v(246)
    assign sha_core_block_next[151] = sha_state_idle ? 1'b0 : n1372;   // sha_top.v(246)
    assign sha_core_block_next[150] = sha_state_idle ? 1'b0 : n1373;   // sha_top.v(246)
    assign sha_core_block_next[149] = sha_state_idle ? 1'b0 : n1374;   // sha_top.v(246)
    assign sha_core_block_next[148] = sha_state_idle ? 1'b0 : n1375;   // sha_top.v(246)
    assign sha_core_block_next[147] = sha_state_idle ? 1'b0 : n1376;   // sha_top.v(246)
    assign sha_core_block_next[146] = sha_state_idle ? 1'b0 : n1377;   // sha_top.v(246)
    assign sha_core_block_next[145] = sha_state_idle ? 1'b0 : n1378;   // sha_top.v(246)
    assign sha_core_block_next[144] = sha_state_idle ? 1'b0 : n1379;   // sha_top.v(246)
    assign sha_core_block_next[143] = sha_state_idle ? 1'b0 : n1380;   // sha_top.v(246)
    assign sha_core_block_next[142] = sha_state_idle ? 1'b0 : n1381;   // sha_top.v(246)
    assign sha_core_block_next[141] = sha_state_idle ? 1'b0 : n1382;   // sha_top.v(246)
    assign sha_core_block_next[140] = sha_state_idle ? 1'b0 : n1383;   // sha_top.v(246)
    assign sha_core_block_next[139] = sha_state_idle ? 1'b0 : n1384;   // sha_top.v(246)
    assign sha_core_block_next[138] = sha_state_idle ? 1'b0 : n1385;   // sha_top.v(246)
    assign sha_core_block_next[137] = sha_state_idle ? 1'b0 : n1386;   // sha_top.v(246)
    assign sha_core_block_next[136] = sha_state_idle ? 1'b0 : n1387;   // sha_top.v(246)
    assign sha_core_block_next[135] = sha_state_idle ? 1'b0 : n1388;   // sha_top.v(246)
    assign sha_core_block_next[134] = sha_state_idle ? 1'b0 : n1389;   // sha_top.v(246)
    assign sha_core_block_next[133] = sha_state_idle ? 1'b0 : n1390;   // sha_top.v(246)
    assign sha_core_block_next[132] = sha_state_idle ? 1'b0 : n1391;   // sha_top.v(246)
    assign sha_core_block_next[131] = sha_state_idle ? 1'b0 : n1392;   // sha_top.v(246)
    assign sha_core_block_next[130] = sha_state_idle ? 1'b0 : n1393;   // sha_top.v(246)
    assign sha_core_block_next[129] = sha_state_idle ? 1'b0 : n1394;   // sha_top.v(246)
    assign sha_core_block_next[128] = sha_state_idle ? 1'b0 : n1395;   // sha_top.v(246)
    assign sha_core_block_next[127] = sha_state_idle ? 1'b0 : n1396;   // sha_top.v(246)
    assign sha_core_block_next[126] = sha_state_idle ? 1'b0 : n1397;   // sha_top.v(246)
    assign sha_core_block_next[125] = sha_state_idle ? 1'b0 : n1398;   // sha_top.v(246)
    assign sha_core_block_next[124] = sha_state_idle ? 1'b0 : n1399;   // sha_top.v(246)
    assign sha_core_block_next[123] = sha_state_idle ? 1'b0 : n1400;   // sha_top.v(246)
    assign sha_core_block_next[122] = sha_state_idle ? 1'b0 : n1401;   // sha_top.v(246)
    assign sha_core_block_next[121] = sha_state_idle ? 1'b0 : n1402;   // sha_top.v(246)
    assign sha_core_block_next[120] = sha_state_idle ? 1'b0 : n1403;   // sha_top.v(246)
    assign sha_core_block_next[119] = sha_state_idle ? 1'b0 : n1404;   // sha_top.v(246)
    assign sha_core_block_next[118] = sha_state_idle ? 1'b0 : n1405;   // sha_top.v(246)
    assign sha_core_block_next[117] = sha_state_idle ? 1'b0 : n1406;   // sha_top.v(246)
    assign sha_core_block_next[116] = sha_state_idle ? 1'b0 : n1407;   // sha_top.v(246)
    assign sha_core_block_next[115] = sha_state_idle ? 1'b0 : n1408;   // sha_top.v(246)
    assign sha_core_block_next[114] = sha_state_idle ? 1'b0 : n1409;   // sha_top.v(246)
    assign sha_core_block_next[113] = sha_state_idle ? 1'b0 : n1410;   // sha_top.v(246)
    assign sha_core_block_next[112] = sha_state_idle ? 1'b0 : n1411;   // sha_top.v(246)
    assign sha_core_block_next[111] = sha_state_idle ? 1'b0 : n1412;   // sha_top.v(246)
    assign sha_core_block_next[110] = sha_state_idle ? 1'b0 : n1413;   // sha_top.v(246)
    assign sha_core_block_next[109] = sha_state_idle ? 1'b0 : n1414;   // sha_top.v(246)
    assign sha_core_block_next[108] = sha_state_idle ? 1'b0 : n1415;   // sha_top.v(246)
    assign sha_core_block_next[107] = sha_state_idle ? 1'b0 : n1416;   // sha_top.v(246)
    assign sha_core_block_next[106] = sha_state_idle ? 1'b0 : n1417;   // sha_top.v(246)
    assign sha_core_block_next[105] = sha_state_idle ? 1'b0 : n1418;   // sha_top.v(246)
    assign sha_core_block_next[104] = sha_state_idle ? 1'b0 : n1419;   // sha_top.v(246)
    assign sha_core_block_next[103] = sha_state_idle ? 1'b0 : n1420;   // sha_top.v(246)
    assign sha_core_block_next[102] = sha_state_idle ? 1'b0 : n1421;   // sha_top.v(246)
    assign sha_core_block_next[101] = sha_state_idle ? 1'b0 : n1422;   // sha_top.v(246)
    assign sha_core_block_next[100] = sha_state_idle ? 1'b0 : n1423;   // sha_top.v(246)
    assign sha_core_block_next[99] = sha_state_idle ? 1'b0 : n1424;   // sha_top.v(246)
    assign sha_core_block_next[98] = sha_state_idle ? 1'b0 : n1425;   // sha_top.v(246)
    assign sha_core_block_next[97] = sha_state_idle ? 1'b0 : n1426;   // sha_top.v(246)
    assign sha_core_block_next[96] = sha_state_idle ? 1'b0 : n1427;   // sha_top.v(246)
    assign sha_core_block_next[95] = sha_state_idle ? 1'b0 : n1428;   // sha_top.v(246)
    assign sha_core_block_next[94] = sha_state_idle ? 1'b0 : n1429;   // sha_top.v(246)
    assign sha_core_block_next[93] = sha_state_idle ? 1'b0 : n1430;   // sha_top.v(246)
    assign sha_core_block_next[92] = sha_state_idle ? 1'b0 : n1431;   // sha_top.v(246)
    assign sha_core_block_next[91] = sha_state_idle ? 1'b0 : n1432;   // sha_top.v(246)
    assign sha_core_block_next[90] = sha_state_idle ? 1'b0 : n1433;   // sha_top.v(246)
    assign sha_core_block_next[89] = sha_state_idle ? 1'b0 : n1434;   // sha_top.v(246)
    assign sha_core_block_next[88] = sha_state_idle ? 1'b0 : n1435;   // sha_top.v(246)
    assign sha_core_block_next[87] = sha_state_idle ? 1'b0 : n1436;   // sha_top.v(246)
    assign sha_core_block_next[86] = sha_state_idle ? 1'b0 : n1437;   // sha_top.v(246)
    assign sha_core_block_next[85] = sha_state_idle ? 1'b0 : n1438;   // sha_top.v(246)
    assign sha_core_block_next[84] = sha_state_idle ? 1'b0 : n1439;   // sha_top.v(246)
    assign sha_core_block_next[83] = sha_state_idle ? 1'b0 : n1440;   // sha_top.v(246)
    assign sha_core_block_next[82] = sha_state_idle ? 1'b0 : n1441;   // sha_top.v(246)
    assign sha_core_block_next[81] = sha_state_idle ? 1'b0 : n1442;   // sha_top.v(246)
    assign sha_core_block_next[80] = sha_state_idle ? 1'b0 : n1443;   // sha_top.v(246)
    assign sha_core_block_next[79] = sha_state_idle ? 1'b0 : n1444;   // sha_top.v(246)
    assign sha_core_block_next[78] = sha_state_idle ? 1'b0 : n1445;   // sha_top.v(246)
    assign sha_core_block_next[77] = sha_state_idle ? 1'b0 : n1446;   // sha_top.v(246)
    assign sha_core_block_next[76] = sha_state_idle ? 1'b0 : n1447;   // sha_top.v(246)
    assign sha_core_block_next[75] = sha_state_idle ? 1'b0 : n1448;   // sha_top.v(246)
    assign sha_core_block_next[74] = sha_state_idle ? 1'b0 : n1449;   // sha_top.v(246)
    assign sha_core_block_next[73] = sha_state_idle ? 1'b0 : n1450;   // sha_top.v(246)
    assign sha_core_block_next[72] = sha_state_idle ? 1'b0 : n1451;   // sha_top.v(246)
    assign sha_core_block_next[71] = sha_state_idle ? 1'b0 : n1452;   // sha_top.v(246)
    assign sha_core_block_next[70] = sha_state_idle ? 1'b0 : n1453;   // sha_top.v(246)
    assign sha_core_block_next[69] = sha_state_idle ? 1'b0 : n1454;   // sha_top.v(246)
    assign sha_core_block_next[68] = sha_state_idle ? 1'b0 : n1455;   // sha_top.v(246)
    assign sha_core_block_next[67] = sha_state_idle ? 1'b0 : n1456;   // sha_top.v(246)
    assign sha_core_block_next[66] = sha_state_idle ? 1'b0 : n1457;   // sha_top.v(246)
    assign sha_core_block_next[65] = sha_state_idle ? 1'b0 : n1458;   // sha_top.v(246)
    assign sha_core_block_next[64] = sha_state_idle ? 1'b0 : n1459;   // sha_top.v(246)
    assign sha_core_block_next[63] = sha_state_idle ? 1'b0 : n1460;   // sha_top.v(246)
    assign sha_core_block_next[62] = sha_state_idle ? 1'b0 : n1461;   // sha_top.v(246)
    assign sha_core_block_next[61] = sha_state_idle ? 1'b0 : n1462;   // sha_top.v(246)
    assign sha_core_block_next[60] = sha_state_idle ? 1'b0 : n1463;   // sha_top.v(246)
    assign sha_core_block_next[59] = sha_state_idle ? 1'b0 : n1464;   // sha_top.v(246)
    assign sha_core_block_next[58] = sha_state_idle ? 1'b0 : n1465;   // sha_top.v(246)
    assign sha_core_block_next[57] = sha_state_idle ? 1'b0 : n1466;   // sha_top.v(246)
    assign sha_core_block_next[56] = sha_state_idle ? 1'b0 : n1467;   // sha_top.v(246)
    assign sha_core_block_next[55] = sha_state_idle ? 1'b0 : n1468;   // sha_top.v(246)
    assign sha_core_block_next[54] = sha_state_idle ? 1'b0 : n1469;   // sha_top.v(246)
    assign sha_core_block_next[53] = sha_state_idle ? 1'b0 : n1470;   // sha_top.v(246)
    assign sha_core_block_next[52] = sha_state_idle ? 1'b0 : n1471;   // sha_top.v(246)
    assign sha_core_block_next[51] = sha_state_idle ? 1'b0 : n1472;   // sha_top.v(246)
    assign sha_core_block_next[50] = sha_state_idle ? 1'b0 : n1473;   // sha_top.v(246)
    assign sha_core_block_next[49] = sha_state_idle ? 1'b0 : n1474;   // sha_top.v(246)
    assign sha_core_block_next[48] = sha_state_idle ? 1'b0 : n1475;   // sha_top.v(246)
    assign sha_core_block_next[47] = sha_state_idle ? 1'b0 : n1476;   // sha_top.v(246)
    assign sha_core_block_next[46] = sha_state_idle ? 1'b0 : n1477;   // sha_top.v(246)
    assign sha_core_block_next[45] = sha_state_idle ? 1'b0 : n1478;   // sha_top.v(246)
    assign sha_core_block_next[44] = sha_state_idle ? 1'b0 : n1479;   // sha_top.v(246)
    assign sha_core_block_next[43] = sha_state_idle ? 1'b0 : n1480;   // sha_top.v(246)
    assign sha_core_block_next[42] = sha_state_idle ? 1'b0 : n1481;   // sha_top.v(246)
    assign sha_core_block_next[41] = sha_state_idle ? 1'b0 : n1482;   // sha_top.v(246)
    assign sha_core_block_next[40] = sha_state_idle ? 1'b0 : n1483;   // sha_top.v(246)
    assign sha_core_block_next[39] = sha_state_idle ? 1'b0 : n1484;   // sha_top.v(246)
    assign sha_core_block_next[38] = sha_state_idle ? 1'b0 : n1485;   // sha_top.v(246)
    assign sha_core_block_next[37] = sha_state_idle ? 1'b0 : n1486;   // sha_top.v(246)
    assign sha_core_block_next[36] = sha_state_idle ? 1'b0 : n1487;   // sha_top.v(246)
    assign sha_core_block_next[35] = sha_state_idle ? 1'b0 : n1488;   // sha_top.v(246)
    assign sha_core_block_next[34] = sha_state_idle ? 1'b0 : n1489;   // sha_top.v(246)
    assign sha_core_block_next[33] = sha_state_idle ? 1'b0 : n1490;   // sha_top.v(246)
    assign sha_core_block_next[32] = sha_state_idle ? 1'b0 : n1491;   // sha_top.v(246)
    assign sha_core_block_next[31] = sha_state_idle ? 1'b0 : n1492;   // sha_top.v(246)
    assign sha_core_block_next[30] = sha_state_idle ? 1'b0 : n1493;   // sha_top.v(246)
    assign sha_core_block_next[29] = sha_state_idle ? 1'b0 : n1494;   // sha_top.v(246)
    assign sha_core_block_next[28] = sha_state_idle ? 1'b0 : n1495;   // sha_top.v(246)
    assign sha_core_block_next[27] = sha_state_idle ? 1'b0 : n1496;   // sha_top.v(246)
    assign sha_core_block_next[26] = sha_state_idle ? 1'b0 : n1497;   // sha_top.v(246)
    assign sha_core_block_next[25] = sha_state_idle ? 1'b0 : n1498;   // sha_top.v(246)
    assign sha_core_block_next[24] = sha_state_idle ? 1'b0 : n1499;   // sha_top.v(246)
    assign sha_core_block_next[23] = sha_state_idle ? 1'b0 : n1500;   // sha_top.v(246)
    assign sha_core_block_next[22] = sha_state_idle ? 1'b0 : n1501;   // sha_top.v(246)
    assign sha_core_block_next[21] = sha_state_idle ? 1'b0 : n1502;   // sha_top.v(246)
    assign sha_core_block_next[20] = sha_state_idle ? 1'b0 : n1503;   // sha_top.v(246)
    assign sha_core_block_next[19] = sha_state_idle ? 1'b0 : n1504;   // sha_top.v(246)
    assign sha_core_block_next[18] = sha_state_idle ? 1'b0 : n1505;   // sha_top.v(246)
    assign sha_core_block_next[17] = sha_state_idle ? 1'b0 : n1506;   // sha_top.v(246)
    assign sha_core_block_next[16] = sha_state_idle ? 1'b0 : n1507;   // sha_top.v(246)
    assign sha_core_block_next[15] = sha_state_idle ? 1'b0 : n1508;   // sha_top.v(246)
    assign sha_core_block_next[14] = sha_state_idle ? 1'b0 : n1509;   // sha_top.v(246)
    assign sha_core_block_next[13] = sha_state_idle ? 1'b0 : n1510;   // sha_top.v(246)
    assign sha_core_block_next[12] = sha_state_idle ? 1'b0 : n1511;   // sha_top.v(246)
    assign sha_core_block_next[11] = sha_state_idle ? 1'b0 : n1512;   // sha_top.v(246)
    assign sha_core_block_next[10] = sha_state_idle ? 1'b0 : n1513;   // sha_top.v(246)
    assign sha_core_block_next[9] = sha_state_idle ? 1'b0 : n1514;   // sha_top.v(246)
    assign sha_core_block_next[8] = sha_state_idle ? 1'b0 : n1515;   // sha_top.v(246)
    assign sha_core_block_next[7] = sha_state_idle ? 1'b0 : n1516;   // sha_top.v(246)
    assign sha_core_block_next[6] = sha_state_idle ? 1'b0 : n1517;   // sha_top.v(246)
    assign sha_core_block_next[5] = sha_state_idle ? 1'b0 : n1518;   // sha_top.v(246)
    assign sha_core_block_next[4] = sha_state_idle ? 1'b0 : n1519;   // sha_top.v(246)
    assign sha_core_block_next[3] = sha_state_idle ? 1'b0 : n1520;   // sha_top.v(246)
    assign sha_core_block_next[2] = sha_state_idle ? 1'b0 : n1521;   // sha_top.v(246)
    assign sha_core_block_next[1] = sha_state_idle ? 1'b0 : n1522;   // sha_top.v(246)
    assign sha_core_block_next[0] = sha_state_idle ? 1'b0 : n1523;   // sha_top.v(246)
    and (write_last_byte_acked, writing_last_byte, xram_ack) ;   // sha_top.v(251)
    assign n2041 = sel_reg_len ? data_out_len[7] : 1'b0;   // sha_top.v(266)
    assign n2042 = sel_reg_len ? data_out_len[6] : 1'b0;   // sha_top.v(266)
    assign n2043 = sel_reg_len ? data_out_len[5] : 1'b0;   // sha_top.v(266)
    assign n2044 = sel_reg_len ? data_out_len[4] : 1'b0;   // sha_top.v(266)
    assign n2045 = sel_reg_len ? data_out_len[3] : 1'b0;   // sha_top.v(266)
    assign n2046 = sel_reg_len ? data_out_len[2] : 1'b0;   // sha_top.v(266)
    assign n2047 = sel_reg_len ? data_out_len[1] : 1'b0;   // sha_top.v(266)
    assign n2048 = sel_reg_len ? data_out_len[0] : 1'b0;   // sha_top.v(266)
    assign n2049 = sel_reg_wr_addr ? data_out_wr_addr[7] : n2041;   // sha_top.v(266)
    assign n2050 = sel_reg_wr_addr ? data_out_wr_addr[6] : n2042;   // sha_top.v(266)
    assign n2051 = sel_reg_wr_addr ? data_out_wr_addr[5] : n2043;   // sha_top.v(266)
    assign n2052 = sel_reg_wr_addr ? data_out_wr_addr[4] : n2044;   // sha_top.v(266)
    assign n2053 = sel_reg_wr_addr ? data_out_wr_addr[3] : n2045;   // sha_top.v(266)
    assign n2054 = sel_reg_wr_addr ? data_out_wr_addr[2] : n2046;   // sha_top.v(266)
    assign n2055 = sel_reg_wr_addr ? data_out_wr_addr[1] : n2047;   // sha_top.v(266)
    assign n2056 = sel_reg_wr_addr ? data_out_wr_addr[0] : n2048;   // sha_top.v(266)
    assign n2057 = sel_reg_rd_addr ? data_out_rd_addr[7] : n2049;   // sha_top.v(266)
    assign n2058 = sel_reg_rd_addr ? data_out_rd_addr[6] : n2050;   // sha_top.v(266)
    assign n2059 = sel_reg_rd_addr ? data_out_rd_addr[5] : n2051;   // sha_top.v(266)
    assign n2060 = sel_reg_rd_addr ? data_out_rd_addr[4] : n2052;   // sha_top.v(266)
    assign n2061 = sel_reg_rd_addr ? data_out_rd_addr[3] : n2053;   // sha_top.v(266)
    assign n2062 = sel_reg_rd_addr ? data_out_rd_addr[2] : n2054;   // sha_top.v(266)
    assign n2063 = sel_reg_rd_addr ? data_out_rd_addr[1] : n2055;   // sha_top.v(266)
    assign n2064 = sel_reg_rd_addr ? data_out_rd_addr[0] : n2056;   // sha_top.v(266)
    assign data_out[7] = sel_reg_state ? 1'b0 : n2057;   // sha_top.v(266)
    assign data_out[6] = sel_reg_state ? 1'b0 : n2058;   // sha_top.v(266)
    assign data_out[5] = sel_reg_state ? 1'b0 : n2059;   // sha_top.v(266)
    assign data_out[4] = sel_reg_state ? 1'b0 : n2060;   // sha_top.v(266)
    assign data_out[3] = sel_reg_state ? 1'b0 : n2061;   // sha_top.v(266)
    assign data_out[2] = sel_reg_state ? sha_state[2] : n2062;   // sha_top.v(266)
    assign data_out[1] = sel_reg_state ? sha_state[1] : n2063;   // sha_top.v(266)
    assign data_out[0] = sel_reg_state ? sha_state[0] : n2064;   // sha_top.v(266)
    reg2byte sha_reg_rd_addr_i (.clk(clk), .rst(rst), .en(sel_reg_rd_addr), 
            .wr(n2073), .addr(addr[0]), .data_in({data_in}), .data_out({data_out_rd_addr}), 
            .reg_out({sha_rdaddr}));   // sha_top.v(270)
    and (n2073, sel_reg_rd_addr, wren) ;   // sha_top.v(274)
    reg2byte sha_reg_wr_addr_i (.clk(clk), .rst(rst), .en(sel_reg_wr_addr), 
            .wr(n2074), .addr(addr[0]), .data_in({data_in}), .data_out({data_out_wr_addr}), 
            .reg_out({sha_wraddr}));   // sha_top.v(283)
    and (n2074, sel_reg_wr_addr, wren) ;   // sha_top.v(287)
    reg2byte sha_reg_len_i (.clk(clk), .rst(rst), .en(sel_reg_len), .wr(n2075), 
            .addr(addr[0]), .data_in({data_in}), .data_out({data_out_len}), 
            .reg_out({sha_len}));   // sha_top.v(296)
    and (n2075, sel_reg_len, wren) ;   // sha_top.v(300)
    not (sha_core_rst_n, rst) ;   // sha_top.v(312)
    and (n2077, sha_state_op1, sha_core_ready_r) ;   // sha_top.v(314)
    nor (n2078, block_counter[15], block_counter[14], block_counter[13], 
        block_counter[12], block_counter[11], block_counter[10], block_counter[9], 
        block_counter[8], block_counter[7], block_counter[6], block_counter[5], 
        block_counter[4], block_counter[3], block_counter[2], block_counter[1], 
        block_counter[0]) ;   // sha_top.v(314)
    and (sha_core_init, n2077, n2078) ;   // sha_top.v(314)
    or (n2081, block_counter[15], block_counter[14], block_counter[13], 
        block_counter[12], block_counter[11], block_counter[10], block_counter[9], 
        block_counter[8], block_counter[7], block_counter[6], block_counter[5], 
        block_counter[4], block_counter[3], block_counter[2], block_counter[1], 
        block_counter[0]) ;   // sha_top.v(316)
    and (sha_core_next, n2077, n2081) ;   // sha_top.v(316)
    assign sha_reg_digest_next[159] = sha_core_digest_valid ? sha_core_digest[159] : sha_reg_digest[159];   // sha_top.v(331)
    assign sha_reg_digest_next[158] = sha_core_digest_valid ? sha_core_digest[158] : sha_reg_digest[158];   // sha_top.v(331)
    assign sha_reg_digest_next[157] = sha_core_digest_valid ? sha_core_digest[157] : sha_reg_digest[157];   // sha_top.v(331)
    assign sha_reg_digest_next[156] = sha_core_digest_valid ? sha_core_digest[156] : sha_reg_digest[156];   // sha_top.v(331)
    assign sha_reg_digest_next[155] = sha_core_digest_valid ? sha_core_digest[155] : sha_reg_digest[155];   // sha_top.v(331)
    assign sha_reg_digest_next[154] = sha_core_digest_valid ? sha_core_digest[154] : sha_reg_digest[154];   // sha_top.v(331)
    assign sha_reg_digest_next[153] = sha_core_digest_valid ? sha_core_digest[153] : sha_reg_digest[153];   // sha_top.v(331)
    assign sha_reg_digest_next[152] = sha_core_digest_valid ? sha_core_digest[152] : sha_reg_digest[152];   // sha_top.v(331)
    assign sha_reg_digest_next[151] = sha_core_digest_valid ? sha_core_digest[151] : sha_reg_digest[151];   // sha_top.v(331)
    assign sha_reg_digest_next[150] = sha_core_digest_valid ? sha_core_digest[150] : sha_reg_digest[150];   // sha_top.v(331)
    assign sha_reg_digest_next[149] = sha_core_digest_valid ? sha_core_digest[149] : sha_reg_digest[149];   // sha_top.v(331)
    assign sha_reg_digest_next[148] = sha_core_digest_valid ? sha_core_digest[148] : sha_reg_digest[148];   // sha_top.v(331)
    assign sha_reg_digest_next[147] = sha_core_digest_valid ? sha_core_digest[147] : sha_reg_digest[147];   // sha_top.v(331)
    assign sha_reg_digest_next[146] = sha_core_digest_valid ? sha_core_digest[146] : sha_reg_digest[146];   // sha_top.v(331)
    assign sha_reg_digest_next[145] = sha_core_digest_valid ? sha_core_digest[145] : sha_reg_digest[145];   // sha_top.v(331)
    assign sha_reg_digest_next[144] = sha_core_digest_valid ? sha_core_digest[144] : sha_reg_digest[144];   // sha_top.v(331)
    assign sha_reg_digest_next[143] = sha_core_digest_valid ? sha_core_digest[143] : sha_reg_digest[143];   // sha_top.v(331)
    assign sha_reg_digest_next[142] = sha_core_digest_valid ? sha_core_digest[142] : sha_reg_digest[142];   // sha_top.v(331)
    assign sha_reg_digest_next[141] = sha_core_digest_valid ? sha_core_digest[141] : sha_reg_digest[141];   // sha_top.v(331)
    assign sha_reg_digest_next[140] = sha_core_digest_valid ? sha_core_digest[140] : sha_reg_digest[140];   // sha_top.v(331)
    assign sha_reg_digest_next[139] = sha_core_digest_valid ? sha_core_digest[139] : sha_reg_digest[139];   // sha_top.v(331)
    assign sha_reg_digest_next[138] = sha_core_digest_valid ? sha_core_digest[138] : sha_reg_digest[138];   // sha_top.v(331)
    assign sha_reg_digest_next[137] = sha_core_digest_valid ? sha_core_digest[137] : sha_reg_digest[137];   // sha_top.v(331)
    assign sha_reg_digest_next[136] = sha_core_digest_valid ? sha_core_digest[136] : sha_reg_digest[136];   // sha_top.v(331)
    assign sha_reg_digest_next[135] = sha_core_digest_valid ? sha_core_digest[135] : sha_reg_digest[135];   // sha_top.v(331)
    assign sha_reg_digest_next[134] = sha_core_digest_valid ? sha_core_digest[134] : sha_reg_digest[134];   // sha_top.v(331)
    assign sha_reg_digest_next[133] = sha_core_digest_valid ? sha_core_digest[133] : sha_reg_digest[133];   // sha_top.v(331)
    assign sha_reg_digest_next[132] = sha_core_digest_valid ? sha_core_digest[132] : sha_reg_digest[132];   // sha_top.v(331)
    assign sha_reg_digest_next[131] = sha_core_digest_valid ? sha_core_digest[131] : sha_reg_digest[131];   // sha_top.v(331)
    assign sha_reg_digest_next[130] = sha_core_digest_valid ? sha_core_digest[130] : sha_reg_digest[130];   // sha_top.v(331)
    assign sha_reg_digest_next[129] = sha_core_digest_valid ? sha_core_digest[129] : sha_reg_digest[129];   // sha_top.v(331)
    assign sha_reg_digest_next[128] = sha_core_digest_valid ? sha_core_digest[128] : sha_reg_digest[128];   // sha_top.v(331)
    assign sha_reg_digest_next[127] = sha_core_digest_valid ? sha_core_digest[127] : sha_reg_digest[127];   // sha_top.v(331)
    assign sha_reg_digest_next[126] = sha_core_digest_valid ? sha_core_digest[126] : sha_reg_digest[126];   // sha_top.v(331)
    assign sha_reg_digest_next[125] = sha_core_digest_valid ? sha_core_digest[125] : sha_reg_digest[125];   // sha_top.v(331)
    assign sha_reg_digest_next[124] = sha_core_digest_valid ? sha_core_digest[124] : sha_reg_digest[124];   // sha_top.v(331)
    assign sha_reg_digest_next[123] = sha_core_digest_valid ? sha_core_digest[123] : sha_reg_digest[123];   // sha_top.v(331)
    assign sha_reg_digest_next[122] = sha_core_digest_valid ? sha_core_digest[122] : sha_reg_digest[122];   // sha_top.v(331)
    assign sha_reg_digest_next[121] = sha_core_digest_valid ? sha_core_digest[121] : sha_reg_digest[121];   // sha_top.v(331)
    assign sha_reg_digest_next[120] = sha_core_digest_valid ? sha_core_digest[120] : sha_reg_digest[120];   // sha_top.v(331)
    assign sha_reg_digest_next[119] = sha_core_digest_valid ? sha_core_digest[119] : sha_reg_digest[119];   // sha_top.v(331)
    assign sha_reg_digest_next[118] = sha_core_digest_valid ? sha_core_digest[118] : sha_reg_digest[118];   // sha_top.v(331)
    assign sha_reg_digest_next[117] = sha_core_digest_valid ? sha_core_digest[117] : sha_reg_digest[117];   // sha_top.v(331)
    assign sha_reg_digest_next[116] = sha_core_digest_valid ? sha_core_digest[116] : sha_reg_digest[116];   // sha_top.v(331)
    assign sha_reg_digest_next[115] = sha_core_digest_valid ? sha_core_digest[115] : sha_reg_digest[115];   // sha_top.v(331)
    assign sha_reg_digest_next[114] = sha_core_digest_valid ? sha_core_digest[114] : sha_reg_digest[114];   // sha_top.v(331)
    assign sha_reg_digest_next[113] = sha_core_digest_valid ? sha_core_digest[113] : sha_reg_digest[113];   // sha_top.v(331)
    assign sha_reg_digest_next[112] = sha_core_digest_valid ? sha_core_digest[112] : sha_reg_digest[112];   // sha_top.v(331)
    assign sha_reg_digest_next[111] = sha_core_digest_valid ? sha_core_digest[111] : sha_reg_digest[111];   // sha_top.v(331)
    assign sha_reg_digest_next[110] = sha_core_digest_valid ? sha_core_digest[110] : sha_reg_digest[110];   // sha_top.v(331)
    assign sha_reg_digest_next[109] = sha_core_digest_valid ? sha_core_digest[109] : sha_reg_digest[109];   // sha_top.v(331)
    assign sha_reg_digest_next[108] = sha_core_digest_valid ? sha_core_digest[108] : sha_reg_digest[108];   // sha_top.v(331)
    assign sha_reg_digest_next[107] = sha_core_digest_valid ? sha_core_digest[107] : sha_reg_digest[107];   // sha_top.v(331)
    assign sha_reg_digest_next[106] = sha_core_digest_valid ? sha_core_digest[106] : sha_reg_digest[106];   // sha_top.v(331)
    assign sha_reg_digest_next[105] = sha_core_digest_valid ? sha_core_digest[105] : sha_reg_digest[105];   // sha_top.v(331)
    assign sha_reg_digest_next[104] = sha_core_digest_valid ? sha_core_digest[104] : sha_reg_digest[104];   // sha_top.v(331)
    assign sha_reg_digest_next[103] = sha_core_digest_valid ? sha_core_digest[103] : sha_reg_digest[103];   // sha_top.v(331)
    assign sha_reg_digest_next[102] = sha_core_digest_valid ? sha_core_digest[102] : sha_reg_digest[102];   // sha_top.v(331)
    assign sha_reg_digest_next[101] = sha_core_digest_valid ? sha_core_digest[101] : sha_reg_digest[101];   // sha_top.v(331)
    assign sha_reg_digest_next[100] = sha_core_digest_valid ? sha_core_digest[100] : sha_reg_digest[100];   // sha_top.v(331)
    assign sha_reg_digest_next[99] = sha_core_digest_valid ? sha_core_digest[99] : sha_reg_digest[99];   // sha_top.v(331)
    assign sha_reg_digest_next[98] = sha_core_digest_valid ? sha_core_digest[98] : sha_reg_digest[98];   // sha_top.v(331)
    assign sha_reg_digest_next[97] = sha_core_digest_valid ? sha_core_digest[97] : sha_reg_digest[97];   // sha_top.v(331)
    assign sha_reg_digest_next[96] = sha_core_digest_valid ? sha_core_digest[96] : sha_reg_digest[96];   // sha_top.v(331)
    assign sha_reg_digest_next[95] = sha_core_digest_valid ? sha_core_digest[95] : sha_reg_digest[95];   // sha_top.v(331)
    assign sha_reg_digest_next[94] = sha_core_digest_valid ? sha_core_digest[94] : sha_reg_digest[94];   // sha_top.v(331)
    assign sha_reg_digest_next[93] = sha_core_digest_valid ? sha_core_digest[93] : sha_reg_digest[93];   // sha_top.v(331)
    assign sha_reg_digest_next[92] = sha_core_digest_valid ? sha_core_digest[92] : sha_reg_digest[92];   // sha_top.v(331)
    assign sha_reg_digest_next[91] = sha_core_digest_valid ? sha_core_digest[91] : sha_reg_digest[91];   // sha_top.v(331)
    assign sha_reg_digest_next[90] = sha_core_digest_valid ? sha_core_digest[90] : sha_reg_digest[90];   // sha_top.v(331)
    assign sha_reg_digest_next[89] = sha_core_digest_valid ? sha_core_digest[89] : sha_reg_digest[89];   // sha_top.v(331)
    assign sha_reg_digest_next[88] = sha_core_digest_valid ? sha_core_digest[88] : sha_reg_digest[88];   // sha_top.v(331)
    assign sha_reg_digest_next[87] = sha_core_digest_valid ? sha_core_digest[87] : sha_reg_digest[87];   // sha_top.v(331)
    assign sha_reg_digest_next[86] = sha_core_digest_valid ? sha_core_digest[86] : sha_reg_digest[86];   // sha_top.v(331)
    assign sha_reg_digest_next[85] = sha_core_digest_valid ? sha_core_digest[85] : sha_reg_digest[85];   // sha_top.v(331)
    assign sha_reg_digest_next[84] = sha_core_digest_valid ? sha_core_digest[84] : sha_reg_digest[84];   // sha_top.v(331)
    assign sha_reg_digest_next[83] = sha_core_digest_valid ? sha_core_digest[83] : sha_reg_digest[83];   // sha_top.v(331)
    assign sha_reg_digest_next[82] = sha_core_digest_valid ? sha_core_digest[82] : sha_reg_digest[82];   // sha_top.v(331)
    assign sha_reg_digest_next[81] = sha_core_digest_valid ? sha_core_digest[81] : sha_reg_digest[81];   // sha_top.v(331)
    assign sha_reg_digest_next[80] = sha_core_digest_valid ? sha_core_digest[80] : sha_reg_digest[80];   // sha_top.v(331)
    assign sha_reg_digest_next[79] = sha_core_digest_valid ? sha_core_digest[79] : sha_reg_digest[79];   // sha_top.v(331)
    assign sha_reg_digest_next[78] = sha_core_digest_valid ? sha_core_digest[78] : sha_reg_digest[78];   // sha_top.v(331)
    assign sha_reg_digest_next[77] = sha_core_digest_valid ? sha_core_digest[77] : sha_reg_digest[77];   // sha_top.v(331)
    assign sha_reg_digest_next[76] = sha_core_digest_valid ? sha_core_digest[76] : sha_reg_digest[76];   // sha_top.v(331)
    assign sha_reg_digest_next[75] = sha_core_digest_valid ? sha_core_digest[75] : sha_reg_digest[75];   // sha_top.v(331)
    assign sha_reg_digest_next[74] = sha_core_digest_valid ? sha_core_digest[74] : sha_reg_digest[74];   // sha_top.v(331)
    assign sha_reg_digest_next[73] = sha_core_digest_valid ? sha_core_digest[73] : sha_reg_digest[73];   // sha_top.v(331)
    assign sha_reg_digest_next[72] = sha_core_digest_valid ? sha_core_digest[72] : sha_reg_digest[72];   // sha_top.v(331)
    assign sha_reg_digest_next[71] = sha_core_digest_valid ? sha_core_digest[71] : sha_reg_digest[71];   // sha_top.v(331)
    assign sha_reg_digest_next[70] = sha_core_digest_valid ? sha_core_digest[70] : sha_reg_digest[70];   // sha_top.v(331)
    assign sha_reg_digest_next[69] = sha_core_digest_valid ? sha_core_digest[69] : sha_reg_digest[69];   // sha_top.v(331)
    assign sha_reg_digest_next[68] = sha_core_digest_valid ? sha_core_digest[68] : sha_reg_digest[68];   // sha_top.v(331)
    assign sha_reg_digest_next[67] = sha_core_digest_valid ? sha_core_digest[67] : sha_reg_digest[67];   // sha_top.v(331)
    assign sha_reg_digest_next[66] = sha_core_digest_valid ? sha_core_digest[66] : sha_reg_digest[66];   // sha_top.v(331)
    assign sha_reg_digest_next[65] = sha_core_digest_valid ? sha_core_digest[65] : sha_reg_digest[65];   // sha_top.v(331)
    assign sha_reg_digest_next[64] = sha_core_digest_valid ? sha_core_digest[64] : sha_reg_digest[64];   // sha_top.v(331)
    assign sha_reg_digest_next[63] = sha_core_digest_valid ? sha_core_digest[63] : sha_reg_digest[63];   // sha_top.v(331)
    assign sha_reg_digest_next[62] = sha_core_digest_valid ? sha_core_digest[62] : sha_reg_digest[62];   // sha_top.v(331)
    assign sha_reg_digest_next[61] = sha_core_digest_valid ? sha_core_digest[61] : sha_reg_digest[61];   // sha_top.v(331)
    assign sha_reg_digest_next[60] = sha_core_digest_valid ? sha_core_digest[60] : sha_reg_digest[60];   // sha_top.v(331)
    assign sha_reg_digest_next[59] = sha_core_digest_valid ? sha_core_digest[59] : sha_reg_digest[59];   // sha_top.v(331)
    assign sha_reg_digest_next[58] = sha_core_digest_valid ? sha_core_digest[58] : sha_reg_digest[58];   // sha_top.v(331)
    assign sha_reg_digest_next[57] = sha_core_digest_valid ? sha_core_digest[57] : sha_reg_digest[57];   // sha_top.v(331)
    assign sha_reg_digest_next[56] = sha_core_digest_valid ? sha_core_digest[56] : sha_reg_digest[56];   // sha_top.v(331)
    assign sha_reg_digest_next[55] = sha_core_digest_valid ? sha_core_digest[55] : sha_reg_digest[55];   // sha_top.v(331)
    assign sha_reg_digest_next[54] = sha_core_digest_valid ? sha_core_digest[54] : sha_reg_digest[54];   // sha_top.v(331)
    assign sha_reg_digest_next[53] = sha_core_digest_valid ? sha_core_digest[53] : sha_reg_digest[53];   // sha_top.v(331)
    assign sha_reg_digest_next[52] = sha_core_digest_valid ? sha_core_digest[52] : sha_reg_digest[52];   // sha_top.v(331)
    assign sha_reg_digest_next[51] = sha_core_digest_valid ? sha_core_digest[51] : sha_reg_digest[51];   // sha_top.v(331)
    assign sha_reg_digest_next[50] = sha_core_digest_valid ? sha_core_digest[50] : sha_reg_digest[50];   // sha_top.v(331)
    assign sha_reg_digest_next[49] = sha_core_digest_valid ? sha_core_digest[49] : sha_reg_digest[49];   // sha_top.v(331)
    assign sha_reg_digest_next[48] = sha_core_digest_valid ? sha_core_digest[48] : sha_reg_digest[48];   // sha_top.v(331)
    assign sha_reg_digest_next[47] = sha_core_digest_valid ? sha_core_digest[47] : sha_reg_digest[47];   // sha_top.v(331)
    assign sha_reg_digest_next[46] = sha_core_digest_valid ? sha_core_digest[46] : sha_reg_digest[46];   // sha_top.v(331)
    assign sha_reg_digest_next[45] = sha_core_digest_valid ? sha_core_digest[45] : sha_reg_digest[45];   // sha_top.v(331)
    assign sha_reg_digest_next[44] = sha_core_digest_valid ? sha_core_digest[44] : sha_reg_digest[44];   // sha_top.v(331)
    assign sha_reg_digest_next[43] = sha_core_digest_valid ? sha_core_digest[43] : sha_reg_digest[43];   // sha_top.v(331)
    assign sha_reg_digest_next[42] = sha_core_digest_valid ? sha_core_digest[42] : sha_reg_digest[42];   // sha_top.v(331)
    assign sha_reg_digest_next[41] = sha_core_digest_valid ? sha_core_digest[41] : sha_reg_digest[41];   // sha_top.v(331)
    assign sha_reg_digest_next[40] = sha_core_digest_valid ? sha_core_digest[40] : sha_reg_digest[40];   // sha_top.v(331)
    assign sha_reg_digest_next[39] = sha_core_digest_valid ? sha_core_digest[39] : sha_reg_digest[39];   // sha_top.v(331)
    assign sha_reg_digest_next[38] = sha_core_digest_valid ? sha_core_digest[38] : sha_reg_digest[38];   // sha_top.v(331)
    assign sha_reg_digest_next[37] = sha_core_digest_valid ? sha_core_digest[37] : sha_reg_digest[37];   // sha_top.v(331)
    assign sha_reg_digest_next[36] = sha_core_digest_valid ? sha_core_digest[36] : sha_reg_digest[36];   // sha_top.v(331)
    assign sha_reg_digest_next[35] = sha_core_digest_valid ? sha_core_digest[35] : sha_reg_digest[35];   // sha_top.v(331)
    assign sha_reg_digest_next[34] = sha_core_digest_valid ? sha_core_digest[34] : sha_reg_digest[34];   // sha_top.v(331)
    assign sha_reg_digest_next[33] = sha_core_digest_valid ? sha_core_digest[33] : sha_reg_digest[33];   // sha_top.v(331)
    assign sha_reg_digest_next[32] = sha_core_digest_valid ? sha_core_digest[32] : sha_reg_digest[32];   // sha_top.v(331)
    assign sha_reg_digest_next[31] = sha_core_digest_valid ? sha_core_digest[31] : sha_reg_digest[31];   // sha_top.v(331)
    assign sha_reg_digest_next[30] = sha_core_digest_valid ? sha_core_digest[30] : sha_reg_digest[30];   // sha_top.v(331)
    assign sha_reg_digest_next[29] = sha_core_digest_valid ? sha_core_digest[29] : sha_reg_digest[29];   // sha_top.v(331)
    assign sha_reg_digest_next[28] = sha_core_digest_valid ? sha_core_digest[28] : sha_reg_digest[28];   // sha_top.v(331)
    assign sha_reg_digest_next[27] = sha_core_digest_valid ? sha_core_digest[27] : sha_reg_digest[27];   // sha_top.v(331)
    assign sha_reg_digest_next[26] = sha_core_digest_valid ? sha_core_digest[26] : sha_reg_digest[26];   // sha_top.v(331)
    assign sha_reg_digest_next[25] = sha_core_digest_valid ? sha_core_digest[25] : sha_reg_digest[25];   // sha_top.v(331)
    assign sha_reg_digest_next[24] = sha_core_digest_valid ? sha_core_digest[24] : sha_reg_digest[24];   // sha_top.v(331)
    assign sha_reg_digest_next[23] = sha_core_digest_valid ? sha_core_digest[23] : sha_reg_digest[23];   // sha_top.v(331)
    assign sha_reg_digest_next[22] = sha_core_digest_valid ? sha_core_digest[22] : sha_reg_digest[22];   // sha_top.v(331)
    assign sha_reg_digest_next[21] = sha_core_digest_valid ? sha_core_digest[21] : sha_reg_digest[21];   // sha_top.v(331)
    assign sha_reg_digest_next[20] = sha_core_digest_valid ? sha_core_digest[20] : sha_reg_digest[20];   // sha_top.v(331)
    assign sha_reg_digest_next[19] = sha_core_digest_valid ? sha_core_digest[19] : sha_reg_digest[19];   // sha_top.v(331)
    assign sha_reg_digest_next[18] = sha_core_digest_valid ? sha_core_digest[18] : sha_reg_digest[18];   // sha_top.v(331)
    assign sha_reg_digest_next[17] = sha_core_digest_valid ? sha_core_digest[17] : sha_reg_digest[17];   // sha_top.v(331)
    assign sha_reg_digest_next[16] = sha_core_digest_valid ? sha_core_digest[16] : sha_reg_digest[16];   // sha_top.v(331)
    assign sha_reg_digest_next[15] = sha_core_digest_valid ? sha_core_digest[15] : sha_reg_digest[15];   // sha_top.v(331)
    assign sha_reg_digest_next[14] = sha_core_digest_valid ? sha_core_digest[14] : sha_reg_digest[14];   // sha_top.v(331)
    assign sha_reg_digest_next[13] = sha_core_digest_valid ? sha_core_digest[13] : sha_reg_digest[13];   // sha_top.v(331)
    assign sha_reg_digest_next[12] = sha_core_digest_valid ? sha_core_digest[12] : sha_reg_digest[12];   // sha_top.v(331)
    assign sha_reg_digest_next[11] = sha_core_digest_valid ? sha_core_digest[11] : sha_reg_digest[11];   // sha_top.v(331)
    assign sha_reg_digest_next[10] = sha_core_digest_valid ? sha_core_digest[10] : sha_reg_digest[10];   // sha_top.v(331)
    assign sha_reg_digest_next[9] = sha_core_digest_valid ? sha_core_digest[9] : sha_reg_digest[9];   // sha_top.v(331)
    assign sha_reg_digest_next[8] = sha_core_digest_valid ? sha_core_digest[8] : sha_reg_digest[8];   // sha_top.v(331)
    assign sha_reg_digest_next[7] = sha_core_digest_valid ? sha_core_digest[7] : sha_reg_digest[7];   // sha_top.v(331)
    assign sha_reg_digest_next[6] = sha_core_digest_valid ? sha_core_digest[6] : sha_reg_digest[6];   // sha_top.v(331)
    assign sha_reg_digest_next[5] = sha_core_digest_valid ? sha_core_digest[5] : sha_reg_digest[5];   // sha_top.v(331)
    assign sha_reg_digest_next[4] = sha_core_digest_valid ? sha_core_digest[4] : sha_reg_digest[4];   // sha_top.v(331)
    assign sha_reg_digest_next[3] = sha_core_digest_valid ? sha_core_digest[3] : sha_reg_digest[3];   // sha_top.v(331)
    assign sha_reg_digest_next[2] = sha_core_digest_valid ? sha_core_digest[2] : sha_reg_digest[2];   // sha_top.v(331)
    assign sha_reg_digest_next[1] = sha_core_digest_valid ? sha_core_digest[1] : sha_reg_digest[1];   // sha_top.v(331)
    assign sha_reg_digest_next[0] = sha_core_digest_valid ? sha_core_digest[0] : sha_reg_digest[0];   // sha_top.v(331)
    VERIFIC_DFFRS i3164 (.d(n2530), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_state[2]));   // sha_top.v(410)
    sha1_core sha1_core_i (.clk(clk), .reset_n(sha_core_rst_n), .init(sha_core_init), 
            .next(sha_core_next), .ready(sha_core_ready), .digest_valid(sha_core_digest_valid), 
            .block({sha_core_block}), .digest({sha_core_digest}));   // sha_top.v(350)
    add_16u_16u add_2216 (.cin(1'b0), .a({sha_rdaddr}), .b({10'b0000000000, 
            byte_counter}), .o({n2250, n2251, n2252, n2253, n2254, 
            n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
            n2263, n2264, n2265}));   // sha_top.v(362)
    add_16u_16u add_2217 (.cin(1'b0), .a({n2250, n2251, n2252, n2253, 
            n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, 
            n2262, n2263, n2264, n2265}), .b({block_counter}), .o({n2267, 
            n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
            n2276, n2277, n2278, n2279, n2280, n2281, n2282}));   // sha_top.v(362)
    add_16u_16u add_2218 (.cin(1'b0), .a({sha_wraddr}), .b({10'b0000000000, 
            byte_counter}), .o({n2284, n2285, n2286, n2287, n2288, 
            n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
            n2297, n2298, n2299}));   // sha_top.v(363)
    assign xram_addr[15] = sha_state_read_data ? n2267 : n2284;   // sha_top.v(363)
    assign xram_addr[14] = sha_state_read_data ? n2268 : n2285;   // sha_top.v(363)
    assign xram_addr[13] = sha_state_read_data ? n2269 : n2286;   // sha_top.v(363)
    assign xram_addr[12] = sha_state_read_data ? n2270 : n2287;   // sha_top.v(363)
    assign xram_addr[11] = sha_state_read_data ? n2271 : n2288;   // sha_top.v(363)
    assign xram_addr[10] = sha_state_read_data ? n2272 : n2289;   // sha_top.v(363)
    assign xram_addr[9] = sha_state_read_data ? n2273 : n2290;   // sha_top.v(363)
    assign xram_addr[8] = sha_state_read_data ? n2274 : n2291;   // sha_top.v(363)
    assign xram_addr[7] = sha_state_read_data ? n2275 : n2292;   // sha_top.v(363)
    assign xram_addr[6] = sha_state_read_data ? n2276 : n2293;   // sha_top.v(363)
    assign xram_addr[5] = sha_state_read_data ? n2277 : n2294;   // sha_top.v(363)
    assign xram_addr[4] = sha_state_read_data ? n2278 : n2295;   // sha_top.v(363)
    assign xram_addr[3] = sha_state_read_data ? n2279 : n2296;   // sha_top.v(363)
    assign xram_addr[2] = sha_state_read_data ? n2280 : n2297;   // sha_top.v(363)
    assign xram_addr[1] = sha_state_read_data ? n2281 : n2298;   // sha_top.v(363)
    assign xram_addr[0] = sha_state_read_data ? n2282 : n2299;   // sha_top.v(363)
    assign n2376 = n994 ? sha_reg_digest[151] : sha_reg_digest[159];   // sha_top.v(384)
    assign n2377 = n994 ? sha_reg_digest[150] : sha_reg_digest[158];   // sha_top.v(384)
    assign n2378 = n994 ? sha_reg_digest[149] : sha_reg_digest[157];   // sha_top.v(384)
    assign n2379 = n994 ? sha_reg_digest[148] : sha_reg_digest[156];   // sha_top.v(384)
    assign n2380 = n994 ? sha_reg_digest[147] : sha_reg_digest[155];   // sha_top.v(384)
    assign n2381 = n994 ? sha_reg_digest[146] : sha_reg_digest[154];   // sha_top.v(384)
    assign n2382 = n994 ? sha_reg_digest[145] : sha_reg_digest[153];   // sha_top.v(384)
    assign n2383 = n994 ? sha_reg_digest[144] : sha_reg_digest[152];   // sha_top.v(384)
    assign n2384 = n984 ? sha_reg_digest[143] : n2376;   // sha_top.v(384)
    assign n2385 = n984 ? sha_reg_digest[142] : n2377;   // sha_top.v(384)
    assign n2386 = n984 ? sha_reg_digest[141] : n2378;   // sha_top.v(384)
    assign n2387 = n984 ? sha_reg_digest[140] : n2379;   // sha_top.v(384)
    assign n2388 = n984 ? sha_reg_digest[139] : n2380;   // sha_top.v(384)
    assign n2389 = n984 ? sha_reg_digest[138] : n2381;   // sha_top.v(384)
    assign n2390 = n984 ? sha_reg_digest[137] : n2382;   // sha_top.v(384)
    assign n2391 = n984 ? sha_reg_digest[136] : n2383;   // sha_top.v(384)
    assign n2392 = n974 ? sha_reg_digest[135] : n2384;   // sha_top.v(384)
    assign n2393 = n974 ? sha_reg_digest[134] : n2385;   // sha_top.v(384)
    assign n2394 = n974 ? sha_reg_digest[133] : n2386;   // sha_top.v(384)
    assign n2395 = n974 ? sha_reg_digest[132] : n2387;   // sha_top.v(384)
    assign n2396 = n974 ? sha_reg_digest[131] : n2388;   // sha_top.v(384)
    assign n2397 = n974 ? sha_reg_digest[130] : n2389;   // sha_top.v(384)
    assign n2398 = n974 ? sha_reg_digest[129] : n2390;   // sha_top.v(384)
    assign n2399 = n974 ? sha_reg_digest[128] : n2391;   // sha_top.v(384)
    assign n2400 = n963 ? sha_reg_digest[127] : n2392;   // sha_top.v(384)
    assign n2401 = n963 ? sha_reg_digest[126] : n2393;   // sha_top.v(384)
    assign n2402 = n963 ? sha_reg_digest[125] : n2394;   // sha_top.v(384)
    assign n2403 = n963 ? sha_reg_digest[124] : n2395;   // sha_top.v(384)
    assign n2404 = n963 ? sha_reg_digest[123] : n2396;   // sha_top.v(384)
    assign n2405 = n963 ? sha_reg_digest[122] : n2397;   // sha_top.v(384)
    assign n2406 = n963 ? sha_reg_digest[121] : n2398;   // sha_top.v(384)
    assign n2407 = n963 ? sha_reg_digest[120] : n2399;   // sha_top.v(384)
    assign n2408 = n953 ? sha_reg_digest[119] : n2400;   // sha_top.v(384)
    assign n2409 = n953 ? sha_reg_digest[118] : n2401;   // sha_top.v(384)
    assign n2410 = n953 ? sha_reg_digest[117] : n2402;   // sha_top.v(384)
    assign n2411 = n953 ? sha_reg_digest[116] : n2403;   // sha_top.v(384)
    assign n2412 = n953 ? sha_reg_digest[115] : n2404;   // sha_top.v(384)
    assign n2413 = n953 ? sha_reg_digest[114] : n2405;   // sha_top.v(384)
    assign n2414 = n953 ? sha_reg_digest[113] : n2406;   // sha_top.v(384)
    assign n2415 = n953 ? sha_reg_digest[112] : n2407;   // sha_top.v(384)
    assign n2416 = n942 ? sha_reg_digest[111] : n2408;   // sha_top.v(384)
    assign n2417 = n942 ? sha_reg_digest[110] : n2409;   // sha_top.v(384)
    assign n2418 = n942 ? sha_reg_digest[109] : n2410;   // sha_top.v(384)
    assign n2419 = n942 ? sha_reg_digest[108] : n2411;   // sha_top.v(384)
    assign n2420 = n942 ? sha_reg_digest[107] : n2412;   // sha_top.v(384)
    assign n2421 = n942 ? sha_reg_digest[106] : n2413;   // sha_top.v(384)
    assign n2422 = n942 ? sha_reg_digest[105] : n2414;   // sha_top.v(384)
    assign n2423 = n942 ? sha_reg_digest[104] : n2415;   // sha_top.v(384)
    assign n2424 = n931 ? sha_reg_digest[103] : n2416;   // sha_top.v(384)
    assign n2425 = n931 ? sha_reg_digest[102] : n2417;   // sha_top.v(384)
    assign n2426 = n931 ? sha_reg_digest[101] : n2418;   // sha_top.v(384)
    assign n2427 = n931 ? sha_reg_digest[100] : n2419;   // sha_top.v(384)
    assign n2428 = n931 ? sha_reg_digest[99] : n2420;   // sha_top.v(384)
    assign n2429 = n931 ? sha_reg_digest[98] : n2421;   // sha_top.v(384)
    assign n2430 = n931 ? sha_reg_digest[97] : n2422;   // sha_top.v(384)
    assign n2431 = n931 ? sha_reg_digest[96] : n2423;   // sha_top.v(384)
    assign n2432 = n919 ? sha_reg_digest[95] : n2424;   // sha_top.v(384)
    assign n2433 = n919 ? sha_reg_digest[94] : n2425;   // sha_top.v(384)
    assign n2434 = n919 ? sha_reg_digest[93] : n2426;   // sha_top.v(384)
    assign n2435 = n919 ? sha_reg_digest[92] : n2427;   // sha_top.v(384)
    assign n2436 = n919 ? sha_reg_digest[91] : n2428;   // sha_top.v(384)
    assign n2437 = n919 ? sha_reg_digest[90] : n2429;   // sha_top.v(384)
    assign n2438 = n919 ? sha_reg_digest[89] : n2430;   // sha_top.v(384)
    assign n2439 = n919 ? sha_reg_digest[88] : n2431;   // sha_top.v(384)
    assign n2440 = n909 ? sha_reg_digest[87] : n2432;   // sha_top.v(384)
    assign n2441 = n909 ? sha_reg_digest[86] : n2433;   // sha_top.v(384)
    assign n2442 = n909 ? sha_reg_digest[85] : n2434;   // sha_top.v(384)
    assign n2443 = n909 ? sha_reg_digest[84] : n2435;   // sha_top.v(384)
    assign n2444 = n909 ? sha_reg_digest[83] : n2436;   // sha_top.v(384)
    assign n2445 = n909 ? sha_reg_digest[82] : n2437;   // sha_top.v(384)
    assign n2446 = n909 ? sha_reg_digest[81] : n2438;   // sha_top.v(384)
    assign n2447 = n909 ? sha_reg_digest[80] : n2439;   // sha_top.v(384)
    assign n2448 = n898 ? sha_reg_digest[79] : n2440;   // sha_top.v(384)
    assign n2449 = n898 ? sha_reg_digest[78] : n2441;   // sha_top.v(384)
    assign n2450 = n898 ? sha_reg_digest[77] : n2442;   // sha_top.v(384)
    assign n2451 = n898 ? sha_reg_digest[76] : n2443;   // sha_top.v(384)
    assign n2452 = n898 ? sha_reg_digest[75] : n2444;   // sha_top.v(384)
    assign n2453 = n898 ? sha_reg_digest[74] : n2445;   // sha_top.v(384)
    assign n2454 = n898 ? sha_reg_digest[73] : n2446;   // sha_top.v(384)
    assign n2455 = n898 ? sha_reg_digest[72] : n2447;   // sha_top.v(384)
    assign n2456 = n887 ? sha_reg_digest[71] : n2448;   // sha_top.v(384)
    assign n2457 = n887 ? sha_reg_digest[70] : n2449;   // sha_top.v(384)
    assign n2458 = n887 ? sha_reg_digest[69] : n2450;   // sha_top.v(384)
    assign n2459 = n887 ? sha_reg_digest[68] : n2451;   // sha_top.v(384)
    assign n2460 = n887 ? sha_reg_digest[67] : n2452;   // sha_top.v(384)
    assign n2461 = n887 ? sha_reg_digest[66] : n2453;   // sha_top.v(384)
    assign n2462 = n887 ? sha_reg_digest[65] : n2454;   // sha_top.v(384)
    assign n2463 = n887 ? sha_reg_digest[64] : n2455;   // sha_top.v(384)
    assign n2464 = n875 ? sha_reg_digest[63] : n2456;   // sha_top.v(384)
    assign n2465 = n875 ? sha_reg_digest[62] : n2457;   // sha_top.v(384)
    assign n2466 = n875 ? sha_reg_digest[61] : n2458;   // sha_top.v(384)
    assign n2467 = n875 ? sha_reg_digest[60] : n2459;   // sha_top.v(384)
    assign n2468 = n875 ? sha_reg_digest[59] : n2460;   // sha_top.v(384)
    assign n2469 = n875 ? sha_reg_digest[58] : n2461;   // sha_top.v(384)
    assign n2470 = n875 ? sha_reg_digest[57] : n2462;   // sha_top.v(384)
    assign n2471 = n875 ? sha_reg_digest[56] : n2463;   // sha_top.v(384)
    assign n2472 = n864 ? sha_reg_digest[55] : n2464;   // sha_top.v(384)
    assign n2473 = n864 ? sha_reg_digest[54] : n2465;   // sha_top.v(384)
    assign n2474 = n864 ? sha_reg_digest[53] : n2466;   // sha_top.v(384)
    assign n2475 = n864 ? sha_reg_digest[52] : n2467;   // sha_top.v(384)
    assign n2476 = n864 ? sha_reg_digest[51] : n2468;   // sha_top.v(384)
    assign n2477 = n864 ? sha_reg_digest[50] : n2469;   // sha_top.v(384)
    assign n2478 = n864 ? sha_reg_digest[49] : n2470;   // sha_top.v(384)
    assign n2479 = n864 ? sha_reg_digest[48] : n2471;   // sha_top.v(384)
    assign n2480 = n852 ? sha_reg_digest[47] : n2472;   // sha_top.v(384)
    assign n2481 = n852 ? sha_reg_digest[46] : n2473;   // sha_top.v(384)
    assign n2482 = n852 ? sha_reg_digest[45] : n2474;   // sha_top.v(384)
    assign n2483 = n852 ? sha_reg_digest[44] : n2475;   // sha_top.v(384)
    assign n2484 = n852 ? sha_reg_digest[43] : n2476;   // sha_top.v(384)
    assign n2485 = n852 ? sha_reg_digest[42] : n2477;   // sha_top.v(384)
    assign n2486 = n852 ? sha_reg_digest[41] : n2478;   // sha_top.v(384)
    assign n2487 = n852 ? sha_reg_digest[40] : n2479;   // sha_top.v(384)
    assign n2488 = n840 ? sha_reg_digest[39] : n2480;   // sha_top.v(384)
    assign n2489 = n840 ? sha_reg_digest[38] : n2481;   // sha_top.v(384)
    assign n2490 = n840 ? sha_reg_digest[37] : n2482;   // sha_top.v(384)
    assign n2491 = n840 ? sha_reg_digest[36] : n2483;   // sha_top.v(384)
    assign n2492 = n840 ? sha_reg_digest[35] : n2484;   // sha_top.v(384)
    assign n2493 = n840 ? sha_reg_digest[34] : n2485;   // sha_top.v(384)
    assign n2494 = n840 ? sha_reg_digest[33] : n2486;   // sha_top.v(384)
    assign n2495 = n840 ? sha_reg_digest[32] : n2487;   // sha_top.v(384)
    assign n2496 = n827 ? sha_reg_digest[31] : n2488;   // sha_top.v(384)
    assign n2497 = n827 ? sha_reg_digest[30] : n2489;   // sha_top.v(384)
    assign n2498 = n827 ? sha_reg_digest[29] : n2490;   // sha_top.v(384)
    assign n2499 = n827 ? sha_reg_digest[28] : n2491;   // sha_top.v(384)
    assign n2500 = n827 ? sha_reg_digest[27] : n2492;   // sha_top.v(384)
    assign n2501 = n827 ? sha_reg_digest[26] : n2493;   // sha_top.v(384)
    assign n2502 = n827 ? sha_reg_digest[25] : n2494;   // sha_top.v(384)
    assign n2503 = n827 ? sha_reg_digest[24] : n2495;   // sha_top.v(384)
    assign n2504 = n817 ? sha_reg_digest[23] : n2496;   // sha_top.v(384)
    assign n2505 = n817 ? sha_reg_digest[22] : n2497;   // sha_top.v(384)
    assign n2506 = n817 ? sha_reg_digest[21] : n2498;   // sha_top.v(384)
    assign n2507 = n817 ? sha_reg_digest[20] : n2499;   // sha_top.v(384)
    assign n2508 = n817 ? sha_reg_digest[19] : n2500;   // sha_top.v(384)
    assign n2509 = n817 ? sha_reg_digest[18] : n2501;   // sha_top.v(384)
    assign n2510 = n817 ? sha_reg_digest[17] : n2502;   // sha_top.v(384)
    assign n2511 = n817 ? sha_reg_digest[16] : n2503;   // sha_top.v(384)
    assign n2512 = n806 ? sha_reg_digest[15] : n2504;   // sha_top.v(384)
    assign n2513 = n806 ? sha_reg_digest[14] : n2505;   // sha_top.v(384)
    assign n2514 = n806 ? sha_reg_digest[13] : n2506;   // sha_top.v(384)
    assign n2515 = n806 ? sha_reg_digest[12] : n2507;   // sha_top.v(384)
    assign n2516 = n806 ? sha_reg_digest[11] : n2508;   // sha_top.v(384)
    assign n2517 = n806 ? sha_reg_digest[10] : n2509;   // sha_top.v(384)
    assign n2518 = n806 ? sha_reg_digest[9] : n2510;   // sha_top.v(384)
    assign n2519 = n806 ? sha_reg_digest[8] : n2511;   // sha_top.v(384)
    assign xram_data_out[7] = writing_last_byte ? sha_reg_digest[7] : n2512;   // sha_top.v(384)
    assign xram_data_out[6] = writing_last_byte ? sha_reg_digest[6] : n2513;   // sha_top.v(384)
    assign xram_data_out[5] = writing_last_byte ? sha_reg_digest[5] : n2514;   // sha_top.v(384)
    assign xram_data_out[4] = writing_last_byte ? sha_reg_digest[4] : n2515;   // sha_top.v(384)
    assign xram_data_out[3] = writing_last_byte ? sha_reg_digest[3] : n2516;   // sha_top.v(384)
    assign xram_data_out[2] = writing_last_byte ? sha_reg_digest[2] : n2517;   // sha_top.v(384)
    assign xram_data_out[1] = writing_last_byte ? sha_reg_digest[1] : n2518;   // sha_top.v(384)
    assign xram_data_out[0] = writing_last_byte ? sha_reg_digest[0] : n2519;   // sha_top.v(384)
    or (xram_stb, sha_state_read_data, xram_wr) ;   // sha_top.v(386)
    assign n2530 = rst ? 1'b0 : sha_state_next[2];   // sha_top.v(409)
    assign n2531 = rst ? 1'b0 : sha_state_next[1];   // sha_top.v(409)
    assign n2532 = rst ? 1'b0 : sha_state_next[0];   // sha_top.v(409)
    assign n2533 = rst ? 1'b0 : byte_counter_next[5];   // sha_top.v(409)
    assign n2534 = rst ? 1'b0 : byte_counter_next[4];   // sha_top.v(409)
    assign n2535 = rst ? 1'b0 : byte_counter_next[3];   // sha_top.v(409)
    assign n2536 = rst ? 1'b0 : byte_counter_next[2];   // sha_top.v(409)
    assign n2537 = rst ? 1'b0 : byte_counter_next[1];   // sha_top.v(409)
    assign n2538 = rst ? 1'b0 : byte_counter_next[0];   // sha_top.v(409)
    assign n2539 = rst ? 1'b0 : sha_core_block_next[511];   // sha_top.v(409)
    assign n2540 = rst ? 1'b0 : sha_core_block_next[510];   // sha_top.v(409)
    assign n2541 = rst ? 1'b0 : sha_core_block_next[509];   // sha_top.v(409)
    assign n2542 = rst ? 1'b0 : sha_core_block_next[508];   // sha_top.v(409)
    assign n2543 = rst ? 1'b0 : sha_core_block_next[507];   // sha_top.v(409)
    assign n2544 = rst ? 1'b0 : sha_core_block_next[506];   // sha_top.v(409)
    assign n2545 = rst ? 1'b0 : sha_core_block_next[505];   // sha_top.v(409)
    assign n2546 = rst ? 1'b0 : sha_core_block_next[504];   // sha_top.v(409)
    assign n2547 = rst ? 1'b0 : sha_core_block_next[503];   // sha_top.v(409)
    assign n2548 = rst ? 1'b0 : sha_core_block_next[502];   // sha_top.v(409)
    assign n2549 = rst ? 1'b0 : sha_core_block_next[501];   // sha_top.v(409)
    assign n2550 = rst ? 1'b0 : sha_core_block_next[500];   // sha_top.v(409)
    assign n2551 = rst ? 1'b0 : sha_core_block_next[499];   // sha_top.v(409)
    assign n2552 = rst ? 1'b0 : sha_core_block_next[498];   // sha_top.v(409)
    assign n2553 = rst ? 1'b0 : sha_core_block_next[497];   // sha_top.v(409)
    assign n2554 = rst ? 1'b0 : sha_core_block_next[496];   // sha_top.v(409)
    assign n2555 = rst ? 1'b0 : sha_core_block_next[495];   // sha_top.v(409)
    assign n2556 = rst ? 1'b0 : sha_core_block_next[494];   // sha_top.v(409)
    assign n2557 = rst ? 1'b0 : sha_core_block_next[493];   // sha_top.v(409)
    assign n2558 = rst ? 1'b0 : sha_core_block_next[492];   // sha_top.v(409)
    assign n2559 = rst ? 1'b0 : sha_core_block_next[491];   // sha_top.v(409)
    assign n2560 = rst ? 1'b0 : sha_core_block_next[490];   // sha_top.v(409)
    assign n2561 = rst ? 1'b0 : sha_core_block_next[489];   // sha_top.v(409)
    assign n2562 = rst ? 1'b0 : sha_core_block_next[488];   // sha_top.v(409)
    assign n2563 = rst ? 1'b0 : sha_core_block_next[487];   // sha_top.v(409)
    assign n2564 = rst ? 1'b0 : sha_core_block_next[486];   // sha_top.v(409)
    assign n2565 = rst ? 1'b0 : sha_core_block_next[485];   // sha_top.v(409)
    assign n2566 = rst ? 1'b0 : sha_core_block_next[484];   // sha_top.v(409)
    assign n2567 = rst ? 1'b0 : sha_core_block_next[483];   // sha_top.v(409)
    assign n2568 = rst ? 1'b0 : sha_core_block_next[482];   // sha_top.v(409)
    assign n2569 = rst ? 1'b0 : sha_core_block_next[481];   // sha_top.v(409)
    assign n2570 = rst ? 1'b0 : sha_core_block_next[480];   // sha_top.v(409)
    assign n2571 = rst ? 1'b0 : sha_core_block_next[479];   // sha_top.v(409)
    assign n2572 = rst ? 1'b0 : sha_core_block_next[478];   // sha_top.v(409)
    assign n2573 = rst ? 1'b0 : sha_core_block_next[477];   // sha_top.v(409)
    assign n2574 = rst ? 1'b0 : sha_core_block_next[476];   // sha_top.v(409)
    assign n2575 = rst ? 1'b0 : sha_core_block_next[475];   // sha_top.v(409)
    assign n2576 = rst ? 1'b0 : sha_core_block_next[474];   // sha_top.v(409)
    assign n2577 = rst ? 1'b0 : sha_core_block_next[473];   // sha_top.v(409)
    assign n2578 = rst ? 1'b0 : sha_core_block_next[472];   // sha_top.v(409)
    assign n2579 = rst ? 1'b0 : sha_core_block_next[471];   // sha_top.v(409)
    assign n2580 = rst ? 1'b0 : sha_core_block_next[470];   // sha_top.v(409)
    assign n2581 = rst ? 1'b0 : sha_core_block_next[469];   // sha_top.v(409)
    assign n2582 = rst ? 1'b0 : sha_core_block_next[468];   // sha_top.v(409)
    assign n2583 = rst ? 1'b0 : sha_core_block_next[467];   // sha_top.v(409)
    assign n2584 = rst ? 1'b0 : sha_core_block_next[466];   // sha_top.v(409)
    assign n2585 = rst ? 1'b0 : sha_core_block_next[465];   // sha_top.v(409)
    assign n2586 = rst ? 1'b0 : sha_core_block_next[464];   // sha_top.v(409)
    assign n2587 = rst ? 1'b0 : sha_core_block_next[463];   // sha_top.v(409)
    assign n2588 = rst ? 1'b0 : sha_core_block_next[462];   // sha_top.v(409)
    assign n2589 = rst ? 1'b0 : sha_core_block_next[461];   // sha_top.v(409)
    assign n2590 = rst ? 1'b0 : sha_core_block_next[460];   // sha_top.v(409)
    assign n2591 = rst ? 1'b0 : sha_core_block_next[459];   // sha_top.v(409)
    assign n2592 = rst ? 1'b0 : sha_core_block_next[458];   // sha_top.v(409)
    assign n2593 = rst ? 1'b0 : sha_core_block_next[457];   // sha_top.v(409)
    assign n2594 = rst ? 1'b0 : sha_core_block_next[456];   // sha_top.v(409)
    assign n2595 = rst ? 1'b0 : sha_core_block_next[455];   // sha_top.v(409)
    assign n2596 = rst ? 1'b0 : sha_core_block_next[454];   // sha_top.v(409)
    assign n2597 = rst ? 1'b0 : sha_core_block_next[453];   // sha_top.v(409)
    assign n2598 = rst ? 1'b0 : sha_core_block_next[452];   // sha_top.v(409)
    assign n2599 = rst ? 1'b0 : sha_core_block_next[451];   // sha_top.v(409)
    assign n2600 = rst ? 1'b0 : sha_core_block_next[450];   // sha_top.v(409)
    assign n2601 = rst ? 1'b0 : sha_core_block_next[449];   // sha_top.v(409)
    assign n2602 = rst ? 1'b0 : sha_core_block_next[448];   // sha_top.v(409)
    assign n2603 = rst ? 1'b0 : sha_core_block_next[447];   // sha_top.v(409)
    assign n2604 = rst ? 1'b0 : sha_core_block_next[446];   // sha_top.v(409)
    assign n2605 = rst ? 1'b0 : sha_core_block_next[445];   // sha_top.v(409)
    assign n2606 = rst ? 1'b0 : sha_core_block_next[444];   // sha_top.v(409)
    assign n2607 = rst ? 1'b0 : sha_core_block_next[443];   // sha_top.v(409)
    assign n2608 = rst ? 1'b0 : sha_core_block_next[442];   // sha_top.v(409)
    assign n2609 = rst ? 1'b0 : sha_core_block_next[441];   // sha_top.v(409)
    assign n2610 = rst ? 1'b0 : sha_core_block_next[440];   // sha_top.v(409)
    assign n2611 = rst ? 1'b0 : sha_core_block_next[439];   // sha_top.v(409)
    assign n2612 = rst ? 1'b0 : sha_core_block_next[438];   // sha_top.v(409)
    assign n2613 = rst ? 1'b0 : sha_core_block_next[437];   // sha_top.v(409)
    assign n2614 = rst ? 1'b0 : sha_core_block_next[436];   // sha_top.v(409)
    assign n2615 = rst ? 1'b0 : sha_core_block_next[435];   // sha_top.v(409)
    assign n2616 = rst ? 1'b0 : sha_core_block_next[434];   // sha_top.v(409)
    assign n2617 = rst ? 1'b0 : sha_core_block_next[433];   // sha_top.v(409)
    assign n2618 = rst ? 1'b0 : sha_core_block_next[432];   // sha_top.v(409)
    assign n2619 = rst ? 1'b0 : sha_core_block_next[431];   // sha_top.v(409)
    assign n2620 = rst ? 1'b0 : sha_core_block_next[430];   // sha_top.v(409)
    assign n2621 = rst ? 1'b0 : sha_core_block_next[429];   // sha_top.v(409)
    assign n2622 = rst ? 1'b0 : sha_core_block_next[428];   // sha_top.v(409)
    assign n2623 = rst ? 1'b0 : sha_core_block_next[427];   // sha_top.v(409)
    assign n2624 = rst ? 1'b0 : sha_core_block_next[426];   // sha_top.v(409)
    assign n2625 = rst ? 1'b0 : sha_core_block_next[425];   // sha_top.v(409)
    assign n2626 = rst ? 1'b0 : sha_core_block_next[424];   // sha_top.v(409)
    assign n2627 = rst ? 1'b0 : sha_core_block_next[423];   // sha_top.v(409)
    assign n2628 = rst ? 1'b0 : sha_core_block_next[422];   // sha_top.v(409)
    assign n2629 = rst ? 1'b0 : sha_core_block_next[421];   // sha_top.v(409)
    assign n2630 = rst ? 1'b0 : sha_core_block_next[420];   // sha_top.v(409)
    assign n2631 = rst ? 1'b0 : sha_core_block_next[419];   // sha_top.v(409)
    assign n2632 = rst ? 1'b0 : sha_core_block_next[418];   // sha_top.v(409)
    assign n2633 = rst ? 1'b0 : sha_core_block_next[417];   // sha_top.v(409)
    assign n2634 = rst ? 1'b0 : sha_core_block_next[416];   // sha_top.v(409)
    assign n2635 = rst ? 1'b0 : sha_core_block_next[415];   // sha_top.v(409)
    assign n2636 = rst ? 1'b0 : sha_core_block_next[414];   // sha_top.v(409)
    assign n2637 = rst ? 1'b0 : sha_core_block_next[413];   // sha_top.v(409)
    assign n2638 = rst ? 1'b0 : sha_core_block_next[412];   // sha_top.v(409)
    assign n2639 = rst ? 1'b0 : sha_core_block_next[411];   // sha_top.v(409)
    assign n2640 = rst ? 1'b0 : sha_core_block_next[410];   // sha_top.v(409)
    assign n2641 = rst ? 1'b0 : sha_core_block_next[409];   // sha_top.v(409)
    assign n2642 = rst ? 1'b0 : sha_core_block_next[408];   // sha_top.v(409)
    assign n2643 = rst ? 1'b0 : sha_core_block_next[407];   // sha_top.v(409)
    assign n2644 = rst ? 1'b0 : sha_core_block_next[406];   // sha_top.v(409)
    assign n2645 = rst ? 1'b0 : sha_core_block_next[405];   // sha_top.v(409)
    assign n2646 = rst ? 1'b0 : sha_core_block_next[404];   // sha_top.v(409)
    assign n2647 = rst ? 1'b0 : sha_core_block_next[403];   // sha_top.v(409)
    assign n2648 = rst ? 1'b0 : sha_core_block_next[402];   // sha_top.v(409)
    assign n2649 = rst ? 1'b0 : sha_core_block_next[401];   // sha_top.v(409)
    assign n2650 = rst ? 1'b0 : sha_core_block_next[400];   // sha_top.v(409)
    assign n2651 = rst ? 1'b0 : sha_core_block_next[399];   // sha_top.v(409)
    assign n2652 = rst ? 1'b0 : sha_core_block_next[398];   // sha_top.v(409)
    assign n2653 = rst ? 1'b0 : sha_core_block_next[397];   // sha_top.v(409)
    assign n2654 = rst ? 1'b0 : sha_core_block_next[396];   // sha_top.v(409)
    assign n2655 = rst ? 1'b0 : sha_core_block_next[395];   // sha_top.v(409)
    assign n2656 = rst ? 1'b0 : sha_core_block_next[394];   // sha_top.v(409)
    assign n2657 = rst ? 1'b0 : sha_core_block_next[393];   // sha_top.v(409)
    assign n2658 = rst ? 1'b0 : sha_core_block_next[392];   // sha_top.v(409)
    assign n2659 = rst ? 1'b0 : sha_core_block_next[391];   // sha_top.v(409)
    assign n2660 = rst ? 1'b0 : sha_core_block_next[390];   // sha_top.v(409)
    assign n2661 = rst ? 1'b0 : sha_core_block_next[389];   // sha_top.v(409)
    assign n2662 = rst ? 1'b0 : sha_core_block_next[388];   // sha_top.v(409)
    assign n2663 = rst ? 1'b0 : sha_core_block_next[387];   // sha_top.v(409)
    assign n2664 = rst ? 1'b0 : sha_core_block_next[386];   // sha_top.v(409)
    assign n2665 = rst ? 1'b0 : sha_core_block_next[385];   // sha_top.v(409)
    assign n2666 = rst ? 1'b0 : sha_core_block_next[384];   // sha_top.v(409)
    assign n2667 = rst ? 1'b0 : sha_core_block_next[383];   // sha_top.v(409)
    assign n2668 = rst ? 1'b0 : sha_core_block_next[382];   // sha_top.v(409)
    assign n2669 = rst ? 1'b0 : sha_core_block_next[381];   // sha_top.v(409)
    assign n2670 = rst ? 1'b0 : sha_core_block_next[380];   // sha_top.v(409)
    assign n2671 = rst ? 1'b0 : sha_core_block_next[379];   // sha_top.v(409)
    assign n2672 = rst ? 1'b0 : sha_core_block_next[378];   // sha_top.v(409)
    assign n2673 = rst ? 1'b0 : sha_core_block_next[377];   // sha_top.v(409)
    assign n2674 = rst ? 1'b0 : sha_core_block_next[376];   // sha_top.v(409)
    assign n2675 = rst ? 1'b0 : sha_core_block_next[375];   // sha_top.v(409)
    assign n2676 = rst ? 1'b0 : sha_core_block_next[374];   // sha_top.v(409)
    assign n2677 = rst ? 1'b0 : sha_core_block_next[373];   // sha_top.v(409)
    assign n2678 = rst ? 1'b0 : sha_core_block_next[372];   // sha_top.v(409)
    assign n2679 = rst ? 1'b0 : sha_core_block_next[371];   // sha_top.v(409)
    assign n2680 = rst ? 1'b0 : sha_core_block_next[370];   // sha_top.v(409)
    assign n2681 = rst ? 1'b0 : sha_core_block_next[369];   // sha_top.v(409)
    assign n2682 = rst ? 1'b0 : sha_core_block_next[368];   // sha_top.v(409)
    assign n2683 = rst ? 1'b0 : sha_core_block_next[367];   // sha_top.v(409)
    assign n2684 = rst ? 1'b0 : sha_core_block_next[366];   // sha_top.v(409)
    assign n2685 = rst ? 1'b0 : sha_core_block_next[365];   // sha_top.v(409)
    assign n2686 = rst ? 1'b0 : sha_core_block_next[364];   // sha_top.v(409)
    assign n2687 = rst ? 1'b0 : sha_core_block_next[363];   // sha_top.v(409)
    assign n2688 = rst ? 1'b0 : sha_core_block_next[362];   // sha_top.v(409)
    assign n2689 = rst ? 1'b0 : sha_core_block_next[361];   // sha_top.v(409)
    assign n2690 = rst ? 1'b0 : sha_core_block_next[360];   // sha_top.v(409)
    assign n2691 = rst ? 1'b0 : sha_core_block_next[359];   // sha_top.v(409)
    assign n2692 = rst ? 1'b0 : sha_core_block_next[358];   // sha_top.v(409)
    assign n2693 = rst ? 1'b0 : sha_core_block_next[357];   // sha_top.v(409)
    assign n2694 = rst ? 1'b0 : sha_core_block_next[356];   // sha_top.v(409)
    assign n2695 = rst ? 1'b0 : sha_core_block_next[355];   // sha_top.v(409)
    assign n2696 = rst ? 1'b0 : sha_core_block_next[354];   // sha_top.v(409)
    assign n2697 = rst ? 1'b0 : sha_core_block_next[353];   // sha_top.v(409)
    assign n2698 = rst ? 1'b0 : sha_core_block_next[352];   // sha_top.v(409)
    assign n2699 = rst ? 1'b0 : sha_core_block_next[351];   // sha_top.v(409)
    assign n2700 = rst ? 1'b0 : sha_core_block_next[350];   // sha_top.v(409)
    assign n2701 = rst ? 1'b0 : sha_core_block_next[349];   // sha_top.v(409)
    assign n2702 = rst ? 1'b0 : sha_core_block_next[348];   // sha_top.v(409)
    assign n2703 = rst ? 1'b0 : sha_core_block_next[347];   // sha_top.v(409)
    assign n2704 = rst ? 1'b0 : sha_core_block_next[346];   // sha_top.v(409)
    assign n2705 = rst ? 1'b0 : sha_core_block_next[345];   // sha_top.v(409)
    assign n2706 = rst ? 1'b0 : sha_core_block_next[344];   // sha_top.v(409)
    assign n2707 = rst ? 1'b0 : sha_core_block_next[343];   // sha_top.v(409)
    assign n2708 = rst ? 1'b0 : sha_core_block_next[342];   // sha_top.v(409)
    assign n2709 = rst ? 1'b0 : sha_core_block_next[341];   // sha_top.v(409)
    assign n2710 = rst ? 1'b0 : sha_core_block_next[340];   // sha_top.v(409)
    assign n2711 = rst ? 1'b0 : sha_core_block_next[339];   // sha_top.v(409)
    assign n2712 = rst ? 1'b0 : sha_core_block_next[338];   // sha_top.v(409)
    assign n2713 = rst ? 1'b0 : sha_core_block_next[337];   // sha_top.v(409)
    assign n2714 = rst ? 1'b0 : sha_core_block_next[336];   // sha_top.v(409)
    assign n2715 = rst ? 1'b0 : sha_core_block_next[335];   // sha_top.v(409)
    assign n2716 = rst ? 1'b0 : sha_core_block_next[334];   // sha_top.v(409)
    assign n2717 = rst ? 1'b0 : sha_core_block_next[333];   // sha_top.v(409)
    assign n2718 = rst ? 1'b0 : sha_core_block_next[332];   // sha_top.v(409)
    assign n2719 = rst ? 1'b0 : sha_core_block_next[331];   // sha_top.v(409)
    assign n2720 = rst ? 1'b0 : sha_core_block_next[330];   // sha_top.v(409)
    assign n2721 = rst ? 1'b0 : sha_core_block_next[329];   // sha_top.v(409)
    assign n2722 = rst ? 1'b0 : sha_core_block_next[328];   // sha_top.v(409)
    assign n2723 = rst ? 1'b0 : sha_core_block_next[327];   // sha_top.v(409)
    assign n2724 = rst ? 1'b0 : sha_core_block_next[326];   // sha_top.v(409)
    assign n2725 = rst ? 1'b0 : sha_core_block_next[325];   // sha_top.v(409)
    assign n2726 = rst ? 1'b0 : sha_core_block_next[324];   // sha_top.v(409)
    assign n2727 = rst ? 1'b0 : sha_core_block_next[323];   // sha_top.v(409)
    assign n2728 = rst ? 1'b0 : sha_core_block_next[322];   // sha_top.v(409)
    assign n2729 = rst ? 1'b0 : sha_core_block_next[321];   // sha_top.v(409)
    assign n2730 = rst ? 1'b0 : sha_core_block_next[320];   // sha_top.v(409)
    assign n2731 = rst ? 1'b0 : sha_core_block_next[319];   // sha_top.v(409)
    assign n2732 = rst ? 1'b0 : sha_core_block_next[318];   // sha_top.v(409)
    assign n2733 = rst ? 1'b0 : sha_core_block_next[317];   // sha_top.v(409)
    assign n2734 = rst ? 1'b0 : sha_core_block_next[316];   // sha_top.v(409)
    assign n2735 = rst ? 1'b0 : sha_core_block_next[315];   // sha_top.v(409)
    assign n2736 = rst ? 1'b0 : sha_core_block_next[314];   // sha_top.v(409)
    assign n2737 = rst ? 1'b0 : sha_core_block_next[313];   // sha_top.v(409)
    assign n2738 = rst ? 1'b0 : sha_core_block_next[312];   // sha_top.v(409)
    assign n2739 = rst ? 1'b0 : sha_core_block_next[311];   // sha_top.v(409)
    assign n2740 = rst ? 1'b0 : sha_core_block_next[310];   // sha_top.v(409)
    assign n2741 = rst ? 1'b0 : sha_core_block_next[309];   // sha_top.v(409)
    assign n2742 = rst ? 1'b0 : sha_core_block_next[308];   // sha_top.v(409)
    assign n2743 = rst ? 1'b0 : sha_core_block_next[307];   // sha_top.v(409)
    assign n2744 = rst ? 1'b0 : sha_core_block_next[306];   // sha_top.v(409)
    assign n2745 = rst ? 1'b0 : sha_core_block_next[305];   // sha_top.v(409)
    assign n2746 = rst ? 1'b0 : sha_core_block_next[304];   // sha_top.v(409)
    assign n2747 = rst ? 1'b0 : sha_core_block_next[303];   // sha_top.v(409)
    assign n2748 = rst ? 1'b0 : sha_core_block_next[302];   // sha_top.v(409)
    assign n2749 = rst ? 1'b0 : sha_core_block_next[301];   // sha_top.v(409)
    assign n2750 = rst ? 1'b0 : sha_core_block_next[300];   // sha_top.v(409)
    assign n2751 = rst ? 1'b0 : sha_core_block_next[299];   // sha_top.v(409)
    assign n2752 = rst ? 1'b0 : sha_core_block_next[298];   // sha_top.v(409)
    assign n2753 = rst ? 1'b0 : sha_core_block_next[297];   // sha_top.v(409)
    assign n2754 = rst ? 1'b0 : sha_core_block_next[296];   // sha_top.v(409)
    assign n2755 = rst ? 1'b0 : sha_core_block_next[295];   // sha_top.v(409)
    assign n2756 = rst ? 1'b0 : sha_core_block_next[294];   // sha_top.v(409)
    assign n2757 = rst ? 1'b0 : sha_core_block_next[293];   // sha_top.v(409)
    assign n2758 = rst ? 1'b0 : sha_core_block_next[292];   // sha_top.v(409)
    assign n2759 = rst ? 1'b0 : sha_core_block_next[291];   // sha_top.v(409)
    assign n2760 = rst ? 1'b0 : sha_core_block_next[290];   // sha_top.v(409)
    assign n2761 = rst ? 1'b0 : sha_core_block_next[289];   // sha_top.v(409)
    assign n2762 = rst ? 1'b0 : sha_core_block_next[288];   // sha_top.v(409)
    assign n2763 = rst ? 1'b0 : sha_core_block_next[287];   // sha_top.v(409)
    assign n2764 = rst ? 1'b0 : sha_core_block_next[286];   // sha_top.v(409)
    assign n2765 = rst ? 1'b0 : sha_core_block_next[285];   // sha_top.v(409)
    assign n2766 = rst ? 1'b0 : sha_core_block_next[284];   // sha_top.v(409)
    assign n2767 = rst ? 1'b0 : sha_core_block_next[283];   // sha_top.v(409)
    assign n2768 = rst ? 1'b0 : sha_core_block_next[282];   // sha_top.v(409)
    assign n2769 = rst ? 1'b0 : sha_core_block_next[281];   // sha_top.v(409)
    assign n2770 = rst ? 1'b0 : sha_core_block_next[280];   // sha_top.v(409)
    assign n2771 = rst ? 1'b0 : sha_core_block_next[279];   // sha_top.v(409)
    assign n2772 = rst ? 1'b0 : sha_core_block_next[278];   // sha_top.v(409)
    assign n2773 = rst ? 1'b0 : sha_core_block_next[277];   // sha_top.v(409)
    assign n2774 = rst ? 1'b0 : sha_core_block_next[276];   // sha_top.v(409)
    assign n2775 = rst ? 1'b0 : sha_core_block_next[275];   // sha_top.v(409)
    assign n2776 = rst ? 1'b0 : sha_core_block_next[274];   // sha_top.v(409)
    assign n2777 = rst ? 1'b0 : sha_core_block_next[273];   // sha_top.v(409)
    assign n2778 = rst ? 1'b0 : sha_core_block_next[272];   // sha_top.v(409)
    assign n2779 = rst ? 1'b0 : sha_core_block_next[271];   // sha_top.v(409)
    assign n2780 = rst ? 1'b0 : sha_core_block_next[270];   // sha_top.v(409)
    assign n2781 = rst ? 1'b0 : sha_core_block_next[269];   // sha_top.v(409)
    assign n2782 = rst ? 1'b0 : sha_core_block_next[268];   // sha_top.v(409)
    assign n2783 = rst ? 1'b0 : sha_core_block_next[267];   // sha_top.v(409)
    assign n2784 = rst ? 1'b0 : sha_core_block_next[266];   // sha_top.v(409)
    assign n2785 = rst ? 1'b0 : sha_core_block_next[265];   // sha_top.v(409)
    assign n2786 = rst ? 1'b0 : sha_core_block_next[264];   // sha_top.v(409)
    assign n2787 = rst ? 1'b0 : sha_core_block_next[263];   // sha_top.v(409)
    assign n2788 = rst ? 1'b0 : sha_core_block_next[262];   // sha_top.v(409)
    assign n2789 = rst ? 1'b0 : sha_core_block_next[261];   // sha_top.v(409)
    assign n2790 = rst ? 1'b0 : sha_core_block_next[260];   // sha_top.v(409)
    assign n2791 = rst ? 1'b0 : sha_core_block_next[259];   // sha_top.v(409)
    assign n2792 = rst ? 1'b0 : sha_core_block_next[258];   // sha_top.v(409)
    assign n2793 = rst ? 1'b0 : sha_core_block_next[257];   // sha_top.v(409)
    assign n2794 = rst ? 1'b0 : sha_core_block_next[256];   // sha_top.v(409)
    assign n2795 = rst ? 1'b0 : sha_core_block_next[255];   // sha_top.v(409)
    assign n2796 = rst ? 1'b0 : sha_core_block_next[254];   // sha_top.v(409)
    assign n2797 = rst ? 1'b0 : sha_core_block_next[253];   // sha_top.v(409)
    assign n2798 = rst ? 1'b0 : sha_core_block_next[252];   // sha_top.v(409)
    assign n2799 = rst ? 1'b0 : sha_core_block_next[251];   // sha_top.v(409)
    assign n2800 = rst ? 1'b0 : sha_core_block_next[250];   // sha_top.v(409)
    assign n2801 = rst ? 1'b0 : sha_core_block_next[249];   // sha_top.v(409)
    assign n2802 = rst ? 1'b0 : sha_core_block_next[248];   // sha_top.v(409)
    assign n2803 = rst ? 1'b0 : sha_core_block_next[247];   // sha_top.v(409)
    assign n2804 = rst ? 1'b0 : sha_core_block_next[246];   // sha_top.v(409)
    assign n2805 = rst ? 1'b0 : sha_core_block_next[245];   // sha_top.v(409)
    assign n2806 = rst ? 1'b0 : sha_core_block_next[244];   // sha_top.v(409)
    assign n2807 = rst ? 1'b0 : sha_core_block_next[243];   // sha_top.v(409)
    assign n2808 = rst ? 1'b0 : sha_core_block_next[242];   // sha_top.v(409)
    assign n2809 = rst ? 1'b0 : sha_core_block_next[241];   // sha_top.v(409)
    assign n2810 = rst ? 1'b0 : sha_core_block_next[240];   // sha_top.v(409)
    assign n2811 = rst ? 1'b0 : sha_core_block_next[239];   // sha_top.v(409)
    assign n2812 = rst ? 1'b0 : sha_core_block_next[238];   // sha_top.v(409)
    assign n2813 = rst ? 1'b0 : sha_core_block_next[237];   // sha_top.v(409)
    assign n2814 = rst ? 1'b0 : sha_core_block_next[236];   // sha_top.v(409)
    assign n2815 = rst ? 1'b0 : sha_core_block_next[235];   // sha_top.v(409)
    assign n2816 = rst ? 1'b0 : sha_core_block_next[234];   // sha_top.v(409)
    assign n2817 = rst ? 1'b0 : sha_core_block_next[233];   // sha_top.v(409)
    assign n2818 = rst ? 1'b0 : sha_core_block_next[232];   // sha_top.v(409)
    assign n2819 = rst ? 1'b0 : sha_core_block_next[231];   // sha_top.v(409)
    assign n2820 = rst ? 1'b0 : sha_core_block_next[230];   // sha_top.v(409)
    assign n2821 = rst ? 1'b0 : sha_core_block_next[229];   // sha_top.v(409)
    assign n2822 = rst ? 1'b0 : sha_core_block_next[228];   // sha_top.v(409)
    assign n2823 = rst ? 1'b0 : sha_core_block_next[227];   // sha_top.v(409)
    assign n2824 = rst ? 1'b0 : sha_core_block_next[226];   // sha_top.v(409)
    assign n2825 = rst ? 1'b0 : sha_core_block_next[225];   // sha_top.v(409)
    assign n2826 = rst ? 1'b0 : sha_core_block_next[224];   // sha_top.v(409)
    assign n2827 = rst ? 1'b0 : sha_core_block_next[223];   // sha_top.v(409)
    assign n2828 = rst ? 1'b0 : sha_core_block_next[222];   // sha_top.v(409)
    assign n2829 = rst ? 1'b0 : sha_core_block_next[221];   // sha_top.v(409)
    assign n2830 = rst ? 1'b0 : sha_core_block_next[220];   // sha_top.v(409)
    assign n2831 = rst ? 1'b0 : sha_core_block_next[219];   // sha_top.v(409)
    assign n2832 = rst ? 1'b0 : sha_core_block_next[218];   // sha_top.v(409)
    assign n2833 = rst ? 1'b0 : sha_core_block_next[217];   // sha_top.v(409)
    assign n2834 = rst ? 1'b0 : sha_core_block_next[216];   // sha_top.v(409)
    assign n2835 = rst ? 1'b0 : sha_core_block_next[215];   // sha_top.v(409)
    assign n2836 = rst ? 1'b0 : sha_core_block_next[214];   // sha_top.v(409)
    assign n2837 = rst ? 1'b0 : sha_core_block_next[213];   // sha_top.v(409)
    assign n2838 = rst ? 1'b0 : sha_core_block_next[212];   // sha_top.v(409)
    assign n2839 = rst ? 1'b0 : sha_core_block_next[211];   // sha_top.v(409)
    assign n2840 = rst ? 1'b0 : sha_core_block_next[210];   // sha_top.v(409)
    assign n2841 = rst ? 1'b0 : sha_core_block_next[209];   // sha_top.v(409)
    assign n2842 = rst ? 1'b0 : sha_core_block_next[208];   // sha_top.v(409)
    assign n2843 = rst ? 1'b0 : sha_core_block_next[207];   // sha_top.v(409)
    assign n2844 = rst ? 1'b0 : sha_core_block_next[206];   // sha_top.v(409)
    assign n2845 = rst ? 1'b0 : sha_core_block_next[205];   // sha_top.v(409)
    assign n2846 = rst ? 1'b0 : sha_core_block_next[204];   // sha_top.v(409)
    assign n2847 = rst ? 1'b0 : sha_core_block_next[203];   // sha_top.v(409)
    assign n2848 = rst ? 1'b0 : sha_core_block_next[202];   // sha_top.v(409)
    assign n2849 = rst ? 1'b0 : sha_core_block_next[201];   // sha_top.v(409)
    assign n2850 = rst ? 1'b0 : sha_core_block_next[200];   // sha_top.v(409)
    assign n2851 = rst ? 1'b0 : sha_core_block_next[199];   // sha_top.v(409)
    assign n2852 = rst ? 1'b0 : sha_core_block_next[198];   // sha_top.v(409)
    assign n2853 = rst ? 1'b0 : sha_core_block_next[197];   // sha_top.v(409)
    assign n2854 = rst ? 1'b0 : sha_core_block_next[196];   // sha_top.v(409)
    assign n2855 = rst ? 1'b0 : sha_core_block_next[195];   // sha_top.v(409)
    assign n2856 = rst ? 1'b0 : sha_core_block_next[194];   // sha_top.v(409)
    assign n2857 = rst ? 1'b0 : sha_core_block_next[193];   // sha_top.v(409)
    assign n2858 = rst ? 1'b0 : sha_core_block_next[192];   // sha_top.v(409)
    assign n2859 = rst ? 1'b0 : sha_core_block_next[191];   // sha_top.v(409)
    assign n2860 = rst ? 1'b0 : sha_core_block_next[190];   // sha_top.v(409)
    assign n2861 = rst ? 1'b0 : sha_core_block_next[189];   // sha_top.v(409)
    assign n2862 = rst ? 1'b0 : sha_core_block_next[188];   // sha_top.v(409)
    assign n2863 = rst ? 1'b0 : sha_core_block_next[187];   // sha_top.v(409)
    assign n2864 = rst ? 1'b0 : sha_core_block_next[186];   // sha_top.v(409)
    assign n2865 = rst ? 1'b0 : sha_core_block_next[185];   // sha_top.v(409)
    assign n2866 = rst ? 1'b0 : sha_core_block_next[184];   // sha_top.v(409)
    assign n2867 = rst ? 1'b0 : sha_core_block_next[183];   // sha_top.v(409)
    assign n2868 = rst ? 1'b0 : sha_core_block_next[182];   // sha_top.v(409)
    assign n2869 = rst ? 1'b0 : sha_core_block_next[181];   // sha_top.v(409)
    assign n2870 = rst ? 1'b0 : sha_core_block_next[180];   // sha_top.v(409)
    assign n2871 = rst ? 1'b0 : sha_core_block_next[179];   // sha_top.v(409)
    assign n2872 = rst ? 1'b0 : sha_core_block_next[178];   // sha_top.v(409)
    assign n2873 = rst ? 1'b0 : sha_core_block_next[177];   // sha_top.v(409)
    assign n2874 = rst ? 1'b0 : sha_core_block_next[176];   // sha_top.v(409)
    assign n2875 = rst ? 1'b0 : sha_core_block_next[175];   // sha_top.v(409)
    assign n2876 = rst ? 1'b0 : sha_core_block_next[174];   // sha_top.v(409)
    assign n2877 = rst ? 1'b0 : sha_core_block_next[173];   // sha_top.v(409)
    assign n2878 = rst ? 1'b0 : sha_core_block_next[172];   // sha_top.v(409)
    assign n2879 = rst ? 1'b0 : sha_core_block_next[171];   // sha_top.v(409)
    assign n2880 = rst ? 1'b0 : sha_core_block_next[170];   // sha_top.v(409)
    assign n2881 = rst ? 1'b0 : sha_core_block_next[169];   // sha_top.v(409)
    assign n2882 = rst ? 1'b0 : sha_core_block_next[168];   // sha_top.v(409)
    assign n2883 = rst ? 1'b0 : sha_core_block_next[167];   // sha_top.v(409)
    assign n2884 = rst ? 1'b0 : sha_core_block_next[166];   // sha_top.v(409)
    assign n2885 = rst ? 1'b0 : sha_core_block_next[165];   // sha_top.v(409)
    assign n2886 = rst ? 1'b0 : sha_core_block_next[164];   // sha_top.v(409)
    assign n2887 = rst ? 1'b0 : sha_core_block_next[163];   // sha_top.v(409)
    assign n2888 = rst ? 1'b0 : sha_core_block_next[162];   // sha_top.v(409)
    assign n2889 = rst ? 1'b0 : sha_core_block_next[161];   // sha_top.v(409)
    assign n2890 = rst ? 1'b0 : sha_core_block_next[160];   // sha_top.v(409)
    assign n2891 = rst ? 1'b0 : sha_core_block_next[159];   // sha_top.v(409)
    assign n2892 = rst ? 1'b0 : sha_core_block_next[158];   // sha_top.v(409)
    assign n2893 = rst ? 1'b0 : sha_core_block_next[157];   // sha_top.v(409)
    assign n2894 = rst ? 1'b0 : sha_core_block_next[156];   // sha_top.v(409)
    assign n2895 = rst ? 1'b0 : sha_core_block_next[155];   // sha_top.v(409)
    assign n2896 = rst ? 1'b0 : sha_core_block_next[154];   // sha_top.v(409)
    assign n2897 = rst ? 1'b0 : sha_core_block_next[153];   // sha_top.v(409)
    assign n2898 = rst ? 1'b0 : sha_core_block_next[152];   // sha_top.v(409)
    assign n2899 = rst ? 1'b0 : sha_core_block_next[151];   // sha_top.v(409)
    assign n2900 = rst ? 1'b0 : sha_core_block_next[150];   // sha_top.v(409)
    assign n2901 = rst ? 1'b0 : sha_core_block_next[149];   // sha_top.v(409)
    assign n2902 = rst ? 1'b0 : sha_core_block_next[148];   // sha_top.v(409)
    assign n2903 = rst ? 1'b0 : sha_core_block_next[147];   // sha_top.v(409)
    assign n2904 = rst ? 1'b0 : sha_core_block_next[146];   // sha_top.v(409)
    assign n2905 = rst ? 1'b0 : sha_core_block_next[145];   // sha_top.v(409)
    assign n2906 = rst ? 1'b0 : sha_core_block_next[144];   // sha_top.v(409)
    assign n2907 = rst ? 1'b0 : sha_core_block_next[143];   // sha_top.v(409)
    assign n2908 = rst ? 1'b0 : sha_core_block_next[142];   // sha_top.v(409)
    assign n2909 = rst ? 1'b0 : sha_core_block_next[141];   // sha_top.v(409)
    assign n2910 = rst ? 1'b0 : sha_core_block_next[140];   // sha_top.v(409)
    assign n2911 = rst ? 1'b0 : sha_core_block_next[139];   // sha_top.v(409)
    assign n2912 = rst ? 1'b0 : sha_core_block_next[138];   // sha_top.v(409)
    assign n2913 = rst ? 1'b0 : sha_core_block_next[137];   // sha_top.v(409)
    assign n2914 = rst ? 1'b0 : sha_core_block_next[136];   // sha_top.v(409)
    assign n2915 = rst ? 1'b0 : sha_core_block_next[135];   // sha_top.v(409)
    assign n2916 = rst ? 1'b0 : sha_core_block_next[134];   // sha_top.v(409)
    assign n2917 = rst ? 1'b0 : sha_core_block_next[133];   // sha_top.v(409)
    assign n2918 = rst ? 1'b0 : sha_core_block_next[132];   // sha_top.v(409)
    assign n2919 = rst ? 1'b0 : sha_core_block_next[131];   // sha_top.v(409)
    assign n2920 = rst ? 1'b0 : sha_core_block_next[130];   // sha_top.v(409)
    assign n2921 = rst ? 1'b0 : sha_core_block_next[129];   // sha_top.v(409)
    assign n2922 = rst ? 1'b0 : sha_core_block_next[128];   // sha_top.v(409)
    assign n2923 = rst ? 1'b0 : sha_core_block_next[127];   // sha_top.v(409)
    assign n2924 = rst ? 1'b0 : sha_core_block_next[126];   // sha_top.v(409)
    assign n2925 = rst ? 1'b0 : sha_core_block_next[125];   // sha_top.v(409)
    assign n2926 = rst ? 1'b0 : sha_core_block_next[124];   // sha_top.v(409)
    assign n2927 = rst ? 1'b0 : sha_core_block_next[123];   // sha_top.v(409)
    assign n2928 = rst ? 1'b0 : sha_core_block_next[122];   // sha_top.v(409)
    assign n2929 = rst ? 1'b0 : sha_core_block_next[121];   // sha_top.v(409)
    assign n2930 = rst ? 1'b0 : sha_core_block_next[120];   // sha_top.v(409)
    assign n2931 = rst ? 1'b0 : sha_core_block_next[119];   // sha_top.v(409)
    assign n2932 = rst ? 1'b0 : sha_core_block_next[118];   // sha_top.v(409)
    assign n2933 = rst ? 1'b0 : sha_core_block_next[117];   // sha_top.v(409)
    assign n2934 = rst ? 1'b0 : sha_core_block_next[116];   // sha_top.v(409)
    assign n2935 = rst ? 1'b0 : sha_core_block_next[115];   // sha_top.v(409)
    assign n2936 = rst ? 1'b0 : sha_core_block_next[114];   // sha_top.v(409)
    assign n2937 = rst ? 1'b0 : sha_core_block_next[113];   // sha_top.v(409)
    assign n2938 = rst ? 1'b0 : sha_core_block_next[112];   // sha_top.v(409)
    assign n2939 = rst ? 1'b0 : sha_core_block_next[111];   // sha_top.v(409)
    assign n2940 = rst ? 1'b0 : sha_core_block_next[110];   // sha_top.v(409)
    assign n2941 = rst ? 1'b0 : sha_core_block_next[109];   // sha_top.v(409)
    assign n2942 = rst ? 1'b0 : sha_core_block_next[108];   // sha_top.v(409)
    assign n2943 = rst ? 1'b0 : sha_core_block_next[107];   // sha_top.v(409)
    assign n2944 = rst ? 1'b0 : sha_core_block_next[106];   // sha_top.v(409)
    assign n2945 = rst ? 1'b0 : sha_core_block_next[105];   // sha_top.v(409)
    assign n2946 = rst ? 1'b0 : sha_core_block_next[104];   // sha_top.v(409)
    assign n2947 = rst ? 1'b0 : sha_core_block_next[103];   // sha_top.v(409)
    assign n2948 = rst ? 1'b0 : sha_core_block_next[102];   // sha_top.v(409)
    assign n2949 = rst ? 1'b0 : sha_core_block_next[101];   // sha_top.v(409)
    assign n2950 = rst ? 1'b0 : sha_core_block_next[100];   // sha_top.v(409)
    assign n2951 = rst ? 1'b0 : sha_core_block_next[99];   // sha_top.v(409)
    assign n2952 = rst ? 1'b0 : sha_core_block_next[98];   // sha_top.v(409)
    assign n2953 = rst ? 1'b0 : sha_core_block_next[97];   // sha_top.v(409)
    assign n2954 = rst ? 1'b0 : sha_core_block_next[96];   // sha_top.v(409)
    assign n2955 = rst ? 1'b0 : sha_core_block_next[95];   // sha_top.v(409)
    assign n2956 = rst ? 1'b0 : sha_core_block_next[94];   // sha_top.v(409)
    assign n2957 = rst ? 1'b0 : sha_core_block_next[93];   // sha_top.v(409)
    assign n2958 = rst ? 1'b0 : sha_core_block_next[92];   // sha_top.v(409)
    assign n2959 = rst ? 1'b0 : sha_core_block_next[91];   // sha_top.v(409)
    assign n2960 = rst ? 1'b0 : sha_core_block_next[90];   // sha_top.v(409)
    assign n2961 = rst ? 1'b0 : sha_core_block_next[89];   // sha_top.v(409)
    assign n2962 = rst ? 1'b0 : sha_core_block_next[88];   // sha_top.v(409)
    assign n2963 = rst ? 1'b0 : sha_core_block_next[87];   // sha_top.v(409)
    assign n2964 = rst ? 1'b0 : sha_core_block_next[86];   // sha_top.v(409)
    assign n2965 = rst ? 1'b0 : sha_core_block_next[85];   // sha_top.v(409)
    assign n2966 = rst ? 1'b0 : sha_core_block_next[84];   // sha_top.v(409)
    assign n2967 = rst ? 1'b0 : sha_core_block_next[83];   // sha_top.v(409)
    assign n2968 = rst ? 1'b0 : sha_core_block_next[82];   // sha_top.v(409)
    assign n2969 = rst ? 1'b0 : sha_core_block_next[81];   // sha_top.v(409)
    assign n2970 = rst ? 1'b0 : sha_core_block_next[80];   // sha_top.v(409)
    assign n2971 = rst ? 1'b0 : sha_core_block_next[79];   // sha_top.v(409)
    assign n2972 = rst ? 1'b0 : sha_core_block_next[78];   // sha_top.v(409)
    assign n2973 = rst ? 1'b0 : sha_core_block_next[77];   // sha_top.v(409)
    assign n2974 = rst ? 1'b0 : sha_core_block_next[76];   // sha_top.v(409)
    assign n2975 = rst ? 1'b0 : sha_core_block_next[75];   // sha_top.v(409)
    assign n2976 = rst ? 1'b0 : sha_core_block_next[74];   // sha_top.v(409)
    assign n2977 = rst ? 1'b0 : sha_core_block_next[73];   // sha_top.v(409)
    assign n2978 = rst ? 1'b0 : sha_core_block_next[72];   // sha_top.v(409)
    assign n2979 = rst ? 1'b0 : sha_core_block_next[71];   // sha_top.v(409)
    assign n2980 = rst ? 1'b0 : sha_core_block_next[70];   // sha_top.v(409)
    assign n2981 = rst ? 1'b0 : sha_core_block_next[69];   // sha_top.v(409)
    assign n2982 = rst ? 1'b0 : sha_core_block_next[68];   // sha_top.v(409)
    assign n2983 = rst ? 1'b0 : sha_core_block_next[67];   // sha_top.v(409)
    assign n2984 = rst ? 1'b0 : sha_core_block_next[66];   // sha_top.v(409)
    assign n2985 = rst ? 1'b0 : sha_core_block_next[65];   // sha_top.v(409)
    assign n2986 = rst ? 1'b0 : sha_core_block_next[64];   // sha_top.v(409)
    assign n2987 = rst ? 1'b0 : sha_core_block_next[63];   // sha_top.v(409)
    assign n2988 = rst ? 1'b0 : sha_core_block_next[62];   // sha_top.v(409)
    assign n2989 = rst ? 1'b0 : sha_core_block_next[61];   // sha_top.v(409)
    assign n2990 = rst ? 1'b0 : sha_core_block_next[60];   // sha_top.v(409)
    assign n2991 = rst ? 1'b0 : sha_core_block_next[59];   // sha_top.v(409)
    assign n2992 = rst ? 1'b0 : sha_core_block_next[58];   // sha_top.v(409)
    assign n2993 = rst ? 1'b0 : sha_core_block_next[57];   // sha_top.v(409)
    assign n2994 = rst ? 1'b0 : sha_core_block_next[56];   // sha_top.v(409)
    assign n2995 = rst ? 1'b0 : sha_core_block_next[55];   // sha_top.v(409)
    assign n2996 = rst ? 1'b0 : sha_core_block_next[54];   // sha_top.v(409)
    assign n2997 = rst ? 1'b0 : sha_core_block_next[53];   // sha_top.v(409)
    assign n2998 = rst ? 1'b0 : sha_core_block_next[52];   // sha_top.v(409)
    assign n2999 = rst ? 1'b0 : sha_core_block_next[51];   // sha_top.v(409)
    assign n3000 = rst ? 1'b0 : sha_core_block_next[50];   // sha_top.v(409)
    assign n3001 = rst ? 1'b0 : sha_core_block_next[49];   // sha_top.v(409)
    assign n3002 = rst ? 1'b0 : sha_core_block_next[48];   // sha_top.v(409)
    assign n3003 = rst ? 1'b0 : sha_core_block_next[47];   // sha_top.v(409)
    assign n3004 = rst ? 1'b0 : sha_core_block_next[46];   // sha_top.v(409)
    assign n3005 = rst ? 1'b0 : sha_core_block_next[45];   // sha_top.v(409)
    assign n3006 = rst ? 1'b0 : sha_core_block_next[44];   // sha_top.v(409)
    assign n3007 = rst ? 1'b0 : sha_core_block_next[43];   // sha_top.v(409)
    assign n3008 = rst ? 1'b0 : sha_core_block_next[42];   // sha_top.v(409)
    assign n3009 = rst ? 1'b0 : sha_core_block_next[41];   // sha_top.v(409)
    assign n3010 = rst ? 1'b0 : sha_core_block_next[40];   // sha_top.v(409)
    assign n3011 = rst ? 1'b0 : sha_core_block_next[39];   // sha_top.v(409)
    assign n3012 = rst ? 1'b0 : sha_core_block_next[38];   // sha_top.v(409)
    assign n3013 = rst ? 1'b0 : sha_core_block_next[37];   // sha_top.v(409)
    assign n3014 = rst ? 1'b0 : sha_core_block_next[36];   // sha_top.v(409)
    assign n3015 = rst ? 1'b0 : sha_core_block_next[35];   // sha_top.v(409)
    assign n3016 = rst ? 1'b0 : sha_core_block_next[34];   // sha_top.v(409)
    assign n3017 = rst ? 1'b0 : sha_core_block_next[33];   // sha_top.v(409)
    assign n3018 = rst ? 1'b0 : sha_core_block_next[32];   // sha_top.v(409)
    assign n3019 = rst ? 1'b0 : sha_core_block_next[31];   // sha_top.v(409)
    assign n3020 = rst ? 1'b0 : sha_core_block_next[30];   // sha_top.v(409)
    assign n3021 = rst ? 1'b0 : sha_core_block_next[29];   // sha_top.v(409)
    assign n3022 = rst ? 1'b0 : sha_core_block_next[28];   // sha_top.v(409)
    assign n3023 = rst ? 1'b0 : sha_core_block_next[27];   // sha_top.v(409)
    assign n3024 = rst ? 1'b0 : sha_core_block_next[26];   // sha_top.v(409)
    assign n3025 = rst ? 1'b0 : sha_core_block_next[25];   // sha_top.v(409)
    assign n3026 = rst ? 1'b0 : sha_core_block_next[24];   // sha_top.v(409)
    assign n3027 = rst ? 1'b0 : sha_core_block_next[23];   // sha_top.v(409)
    assign n3028 = rst ? 1'b0 : sha_core_block_next[22];   // sha_top.v(409)
    assign n3029 = rst ? 1'b0 : sha_core_block_next[21];   // sha_top.v(409)
    assign n3030 = rst ? 1'b0 : sha_core_block_next[20];   // sha_top.v(409)
    assign n3031 = rst ? 1'b0 : sha_core_block_next[19];   // sha_top.v(409)
    assign n3032 = rst ? 1'b0 : sha_core_block_next[18];   // sha_top.v(409)
    assign n3033 = rst ? 1'b0 : sha_core_block_next[17];   // sha_top.v(409)
    assign n3034 = rst ? 1'b0 : sha_core_block_next[16];   // sha_top.v(409)
    assign n3035 = rst ? 1'b0 : sha_core_block_next[15];   // sha_top.v(409)
    assign n3036 = rst ? 1'b0 : sha_core_block_next[14];   // sha_top.v(409)
    assign n3037 = rst ? 1'b0 : sha_core_block_next[13];   // sha_top.v(409)
    assign n3038 = rst ? 1'b0 : sha_core_block_next[12];   // sha_top.v(409)
    assign n3039 = rst ? 1'b0 : sha_core_block_next[11];   // sha_top.v(409)
    assign n3040 = rst ? 1'b0 : sha_core_block_next[10];   // sha_top.v(409)
    assign n3041 = rst ? 1'b0 : sha_core_block_next[9];   // sha_top.v(409)
    assign n3042 = rst ? 1'b0 : sha_core_block_next[8];   // sha_top.v(409)
    assign n3043 = rst ? 1'b0 : sha_core_block_next[7];   // sha_top.v(409)
    assign n3044 = rst ? 1'b0 : sha_core_block_next[6];   // sha_top.v(409)
    assign n3045 = rst ? 1'b0 : sha_core_block_next[5];   // sha_top.v(409)
    assign n3046 = rst ? 1'b0 : sha_core_block_next[4];   // sha_top.v(409)
    assign n3047 = rst ? 1'b0 : sha_core_block_next[3];   // sha_top.v(409)
    assign n3048 = rst ? 1'b0 : sha_core_block_next[2];   // sha_top.v(409)
    assign n3049 = rst ? 1'b0 : sha_core_block_next[1];   // sha_top.v(409)
    assign n3050 = rst ? 1'b0 : sha_core_block_next[0];   // sha_top.v(409)
    assign n3051 = rst ? 1'b0 : bytes_read_next[15];   // sha_top.v(409)
    assign n3052 = rst ? 1'b0 : bytes_read_next[14];   // sha_top.v(409)
    assign n3053 = rst ? 1'b0 : bytes_read_next[13];   // sha_top.v(409)
    assign n3054 = rst ? 1'b0 : bytes_read_next[12];   // sha_top.v(409)
    assign n3055 = rst ? 1'b0 : bytes_read_next[11];   // sha_top.v(409)
    assign n3056 = rst ? 1'b0 : bytes_read_next[10];   // sha_top.v(409)
    assign n3057 = rst ? 1'b0 : bytes_read_next[9];   // sha_top.v(409)
    assign n3058 = rst ? 1'b0 : bytes_read_next[8];   // sha_top.v(409)
    assign n3059 = rst ? 1'b0 : bytes_read_next[7];   // sha_top.v(409)
    assign n3060 = rst ? 1'b0 : bytes_read_next[6];   // sha_top.v(409)
    assign n3061 = rst ? 1'b0 : bytes_read_next[5];   // sha_top.v(409)
    assign n3062 = rst ? 1'b0 : bytes_read_next[4];   // sha_top.v(409)
    assign n3063 = rst ? 1'b0 : bytes_read_next[3];   // sha_top.v(409)
    assign n3064 = rst ? 1'b0 : bytes_read_next[2];   // sha_top.v(409)
    assign n3065 = rst ? 1'b0 : bytes_read_next[1];   // sha_top.v(409)
    assign n3066 = rst ? 1'b0 : bytes_read_next[0];   // sha_top.v(409)
    assign n3067 = rst ? 1'b0 : block_counter_next[15];   // sha_top.v(409)
    assign n3068 = rst ? 1'b0 : block_counter_next[14];   // sha_top.v(409)
    assign n3069 = rst ? 1'b0 : block_counter_next[13];   // sha_top.v(409)
    assign n3070 = rst ? 1'b0 : block_counter_next[12];   // sha_top.v(409)
    assign n3071 = rst ? 1'b0 : block_counter_next[11];   // sha_top.v(409)
    assign n3072 = rst ? 1'b0 : block_counter_next[10];   // sha_top.v(409)
    assign n3073 = rst ? 1'b0 : block_counter_next[9];   // sha_top.v(409)
    assign n3074 = rst ? 1'b0 : block_counter_next[8];   // sha_top.v(409)
    assign n3075 = rst ? 1'b0 : block_counter_next[7];   // sha_top.v(409)
    assign n3076 = rst ? 1'b0 : block_counter_next[6];   // sha_top.v(409)
    assign n3077 = rst ? 1'b0 : block_counter_next[5];   // sha_top.v(409)
    assign n3078 = rst ? 1'b0 : block_counter_next[4];   // sha_top.v(409)
    assign n3079 = rst ? 1'b0 : block_counter_next[3];   // sha_top.v(409)
    assign n3080 = rst ? 1'b0 : block_counter_next[2];   // sha_top.v(409)
    assign n3081 = rst ? 1'b0 : block_counter_next[1];   // sha_top.v(409)
    assign n3082 = rst ? 1'b0 : block_counter_next[0];   // sha_top.v(409)
    assign n3083 = rst ? 1'b0 : sha_reg_digest_next[159];   // sha_top.v(409)
    assign n3084 = rst ? 1'b0 : sha_reg_digest_next[158];   // sha_top.v(409)
    assign n3085 = rst ? 1'b0 : sha_reg_digest_next[157];   // sha_top.v(409)
    assign n3086 = rst ? 1'b0 : sha_reg_digest_next[156];   // sha_top.v(409)
    assign n3087 = rst ? 1'b0 : sha_reg_digest_next[155];   // sha_top.v(409)
    assign n3088 = rst ? 1'b0 : sha_reg_digest_next[154];   // sha_top.v(409)
    assign n3089 = rst ? 1'b0 : sha_reg_digest_next[153];   // sha_top.v(409)
    assign n3090 = rst ? 1'b0 : sha_reg_digest_next[152];   // sha_top.v(409)
    assign n3091 = rst ? 1'b0 : sha_reg_digest_next[151];   // sha_top.v(409)
    assign n3092 = rst ? 1'b0 : sha_reg_digest_next[150];   // sha_top.v(409)
    assign n3093 = rst ? 1'b0 : sha_reg_digest_next[149];   // sha_top.v(409)
    assign n3094 = rst ? 1'b0 : sha_reg_digest_next[148];   // sha_top.v(409)
    assign n3095 = rst ? 1'b0 : sha_reg_digest_next[147];   // sha_top.v(409)
    assign n3096 = rst ? 1'b0 : sha_reg_digest_next[146];   // sha_top.v(409)
    assign n3097 = rst ? 1'b0 : sha_reg_digest_next[145];   // sha_top.v(409)
    assign n3098 = rst ? 1'b0 : sha_reg_digest_next[144];   // sha_top.v(409)
    assign n3099 = rst ? 1'b0 : sha_reg_digest_next[143];   // sha_top.v(409)
    assign n3100 = rst ? 1'b0 : sha_reg_digest_next[142];   // sha_top.v(409)
    assign n3101 = rst ? 1'b0 : sha_reg_digest_next[141];   // sha_top.v(409)
    assign n3102 = rst ? 1'b0 : sha_reg_digest_next[140];   // sha_top.v(409)
    assign n3103 = rst ? 1'b0 : sha_reg_digest_next[139];   // sha_top.v(409)
    assign n3104 = rst ? 1'b0 : sha_reg_digest_next[138];   // sha_top.v(409)
    assign n3105 = rst ? 1'b0 : sha_reg_digest_next[137];   // sha_top.v(409)
    assign n3106 = rst ? 1'b0 : sha_reg_digest_next[136];   // sha_top.v(409)
    assign n3107 = rst ? 1'b0 : sha_reg_digest_next[135];   // sha_top.v(409)
    assign n3108 = rst ? 1'b0 : sha_reg_digest_next[134];   // sha_top.v(409)
    assign n3109 = rst ? 1'b0 : sha_reg_digest_next[133];   // sha_top.v(409)
    assign n3110 = rst ? 1'b0 : sha_reg_digest_next[132];   // sha_top.v(409)
    assign n3111 = rst ? 1'b0 : sha_reg_digest_next[131];   // sha_top.v(409)
    assign n3112 = rst ? 1'b0 : sha_reg_digest_next[130];   // sha_top.v(409)
    assign n3113 = rst ? 1'b0 : sha_reg_digest_next[129];   // sha_top.v(409)
    assign n3114 = rst ? 1'b0 : sha_reg_digest_next[128];   // sha_top.v(409)
    assign n3115 = rst ? 1'b0 : sha_reg_digest_next[127];   // sha_top.v(409)
    assign n3116 = rst ? 1'b0 : sha_reg_digest_next[126];   // sha_top.v(409)
    assign n3117 = rst ? 1'b0 : sha_reg_digest_next[125];   // sha_top.v(409)
    assign n3118 = rst ? 1'b0 : sha_reg_digest_next[124];   // sha_top.v(409)
    assign n3119 = rst ? 1'b0 : sha_reg_digest_next[123];   // sha_top.v(409)
    assign n3120 = rst ? 1'b0 : sha_reg_digest_next[122];   // sha_top.v(409)
    assign n3121 = rst ? 1'b0 : sha_reg_digest_next[121];   // sha_top.v(409)
    assign n3122 = rst ? 1'b0 : sha_reg_digest_next[120];   // sha_top.v(409)
    assign n3123 = rst ? 1'b0 : sha_reg_digest_next[119];   // sha_top.v(409)
    assign n3124 = rst ? 1'b0 : sha_reg_digest_next[118];   // sha_top.v(409)
    assign n3125 = rst ? 1'b0 : sha_reg_digest_next[117];   // sha_top.v(409)
    assign n3126 = rst ? 1'b0 : sha_reg_digest_next[116];   // sha_top.v(409)
    assign n3127 = rst ? 1'b0 : sha_reg_digest_next[115];   // sha_top.v(409)
    assign n3128 = rst ? 1'b0 : sha_reg_digest_next[114];   // sha_top.v(409)
    assign n3129 = rst ? 1'b0 : sha_reg_digest_next[113];   // sha_top.v(409)
    assign n3130 = rst ? 1'b0 : sha_reg_digest_next[112];   // sha_top.v(409)
    assign n3131 = rst ? 1'b0 : sha_reg_digest_next[111];   // sha_top.v(409)
    assign n3132 = rst ? 1'b0 : sha_reg_digest_next[110];   // sha_top.v(409)
    assign n3133 = rst ? 1'b0 : sha_reg_digest_next[109];   // sha_top.v(409)
    assign n3134 = rst ? 1'b0 : sha_reg_digest_next[108];   // sha_top.v(409)
    assign n3135 = rst ? 1'b0 : sha_reg_digest_next[107];   // sha_top.v(409)
    assign n3136 = rst ? 1'b0 : sha_reg_digest_next[106];   // sha_top.v(409)
    assign n3137 = rst ? 1'b0 : sha_reg_digest_next[105];   // sha_top.v(409)
    assign n3138 = rst ? 1'b0 : sha_reg_digest_next[104];   // sha_top.v(409)
    assign n3139 = rst ? 1'b0 : sha_reg_digest_next[103];   // sha_top.v(409)
    assign n3140 = rst ? 1'b0 : sha_reg_digest_next[102];   // sha_top.v(409)
    assign n3141 = rst ? 1'b0 : sha_reg_digest_next[101];   // sha_top.v(409)
    assign n3142 = rst ? 1'b0 : sha_reg_digest_next[100];   // sha_top.v(409)
    assign n3143 = rst ? 1'b0 : sha_reg_digest_next[99];   // sha_top.v(409)
    assign n3144 = rst ? 1'b0 : sha_reg_digest_next[98];   // sha_top.v(409)
    assign n3145 = rst ? 1'b0 : sha_reg_digest_next[97];   // sha_top.v(409)
    assign n3146 = rst ? 1'b0 : sha_reg_digest_next[96];   // sha_top.v(409)
    assign n3147 = rst ? 1'b0 : sha_reg_digest_next[95];   // sha_top.v(409)
    assign n3148 = rst ? 1'b0 : sha_reg_digest_next[94];   // sha_top.v(409)
    assign n3149 = rst ? 1'b0 : sha_reg_digest_next[93];   // sha_top.v(409)
    assign n3150 = rst ? 1'b0 : sha_reg_digest_next[92];   // sha_top.v(409)
    assign n3151 = rst ? 1'b0 : sha_reg_digest_next[91];   // sha_top.v(409)
    assign n3152 = rst ? 1'b0 : sha_reg_digest_next[90];   // sha_top.v(409)
    assign n3153 = rst ? 1'b0 : sha_reg_digest_next[89];   // sha_top.v(409)
    assign n3154 = rst ? 1'b0 : sha_reg_digest_next[88];   // sha_top.v(409)
    assign n3155 = rst ? 1'b0 : sha_reg_digest_next[87];   // sha_top.v(409)
    assign n3156 = rst ? 1'b0 : sha_reg_digest_next[86];   // sha_top.v(409)
    assign n3157 = rst ? 1'b0 : sha_reg_digest_next[85];   // sha_top.v(409)
    assign n3158 = rst ? 1'b0 : sha_reg_digest_next[84];   // sha_top.v(409)
    assign n3159 = rst ? 1'b0 : sha_reg_digest_next[83];   // sha_top.v(409)
    assign n3160 = rst ? 1'b0 : sha_reg_digest_next[82];   // sha_top.v(409)
    assign n3161 = rst ? 1'b0 : sha_reg_digest_next[81];   // sha_top.v(409)
    assign n3162 = rst ? 1'b0 : sha_reg_digest_next[80];   // sha_top.v(409)
    assign n3163 = rst ? 1'b0 : sha_reg_digest_next[79];   // sha_top.v(409)
    assign n3164 = rst ? 1'b0 : sha_reg_digest_next[78];   // sha_top.v(409)
    assign n3165 = rst ? 1'b0 : sha_reg_digest_next[77];   // sha_top.v(409)
    assign n3166 = rst ? 1'b0 : sha_reg_digest_next[76];   // sha_top.v(409)
    assign n3167 = rst ? 1'b0 : sha_reg_digest_next[75];   // sha_top.v(409)
    assign n3168 = rst ? 1'b0 : sha_reg_digest_next[74];   // sha_top.v(409)
    assign n3169 = rst ? 1'b0 : sha_reg_digest_next[73];   // sha_top.v(409)
    assign n3170 = rst ? 1'b0 : sha_reg_digest_next[72];   // sha_top.v(409)
    assign n3171 = rst ? 1'b0 : sha_reg_digest_next[71];   // sha_top.v(409)
    assign n3172 = rst ? 1'b0 : sha_reg_digest_next[70];   // sha_top.v(409)
    assign n3173 = rst ? 1'b0 : sha_reg_digest_next[69];   // sha_top.v(409)
    assign n3174 = rst ? 1'b0 : sha_reg_digest_next[68];   // sha_top.v(409)
    assign n3175 = rst ? 1'b0 : sha_reg_digest_next[67];   // sha_top.v(409)
    assign n3176 = rst ? 1'b0 : sha_reg_digest_next[66];   // sha_top.v(409)
    assign n3177 = rst ? 1'b0 : sha_reg_digest_next[65];   // sha_top.v(409)
    assign n3178 = rst ? 1'b0 : sha_reg_digest_next[64];   // sha_top.v(409)
    assign n3179 = rst ? 1'b0 : sha_reg_digest_next[63];   // sha_top.v(409)
    assign n3180 = rst ? 1'b0 : sha_reg_digest_next[62];   // sha_top.v(409)
    assign n3181 = rst ? 1'b0 : sha_reg_digest_next[61];   // sha_top.v(409)
    assign n3182 = rst ? 1'b0 : sha_reg_digest_next[60];   // sha_top.v(409)
    assign n3183 = rst ? 1'b0 : sha_reg_digest_next[59];   // sha_top.v(409)
    assign n3184 = rst ? 1'b0 : sha_reg_digest_next[58];   // sha_top.v(409)
    assign n3185 = rst ? 1'b0 : sha_reg_digest_next[57];   // sha_top.v(409)
    assign n3186 = rst ? 1'b0 : sha_reg_digest_next[56];   // sha_top.v(409)
    assign n3187 = rst ? 1'b0 : sha_reg_digest_next[55];   // sha_top.v(409)
    assign n3188 = rst ? 1'b0 : sha_reg_digest_next[54];   // sha_top.v(409)
    assign n3189 = rst ? 1'b0 : sha_reg_digest_next[53];   // sha_top.v(409)
    assign n3190 = rst ? 1'b0 : sha_reg_digest_next[52];   // sha_top.v(409)
    assign n3191 = rst ? 1'b0 : sha_reg_digest_next[51];   // sha_top.v(409)
    assign n3192 = rst ? 1'b0 : sha_reg_digest_next[50];   // sha_top.v(409)
    assign n3193 = rst ? 1'b0 : sha_reg_digest_next[49];   // sha_top.v(409)
    assign n3194 = rst ? 1'b0 : sha_reg_digest_next[48];   // sha_top.v(409)
    assign n3195 = rst ? 1'b0 : sha_reg_digest_next[47];   // sha_top.v(409)
    assign n3196 = rst ? 1'b0 : sha_reg_digest_next[46];   // sha_top.v(409)
    assign n3197 = rst ? 1'b0 : sha_reg_digest_next[45];   // sha_top.v(409)
    assign n3198 = rst ? 1'b0 : sha_reg_digest_next[44];   // sha_top.v(409)
    assign n3199 = rst ? 1'b0 : sha_reg_digest_next[43];   // sha_top.v(409)
    assign n3200 = rst ? 1'b0 : sha_reg_digest_next[42];   // sha_top.v(409)
    assign n3201 = rst ? 1'b0 : sha_reg_digest_next[41];   // sha_top.v(409)
    assign n3202 = rst ? 1'b0 : sha_reg_digest_next[40];   // sha_top.v(409)
    assign n3203 = rst ? 1'b0 : sha_reg_digest_next[39];   // sha_top.v(409)
    assign n3204 = rst ? 1'b0 : sha_reg_digest_next[38];   // sha_top.v(409)
    assign n3205 = rst ? 1'b0 : sha_reg_digest_next[37];   // sha_top.v(409)
    assign n3206 = rst ? 1'b0 : sha_reg_digest_next[36];   // sha_top.v(409)
    assign n3207 = rst ? 1'b0 : sha_reg_digest_next[35];   // sha_top.v(409)
    assign n3208 = rst ? 1'b0 : sha_reg_digest_next[34];   // sha_top.v(409)
    assign n3209 = rst ? 1'b0 : sha_reg_digest_next[33];   // sha_top.v(409)
    assign n3210 = rst ? 1'b0 : sha_reg_digest_next[32];   // sha_top.v(409)
    assign n3211 = rst ? 1'b0 : sha_reg_digest_next[31];   // sha_top.v(409)
    assign n3212 = rst ? 1'b0 : sha_reg_digest_next[30];   // sha_top.v(409)
    assign n3213 = rst ? 1'b0 : sha_reg_digest_next[29];   // sha_top.v(409)
    assign n3214 = rst ? 1'b0 : sha_reg_digest_next[28];   // sha_top.v(409)
    assign n3215 = rst ? 1'b0 : sha_reg_digest_next[27];   // sha_top.v(409)
    assign n3216 = rst ? 1'b0 : sha_reg_digest_next[26];   // sha_top.v(409)
    assign n3217 = rst ? 1'b0 : sha_reg_digest_next[25];   // sha_top.v(409)
    assign n3218 = rst ? 1'b0 : sha_reg_digest_next[24];   // sha_top.v(409)
    assign n3219 = rst ? 1'b0 : sha_reg_digest_next[23];   // sha_top.v(409)
    assign n3220 = rst ? 1'b0 : sha_reg_digest_next[22];   // sha_top.v(409)
    assign n3221 = rst ? 1'b0 : sha_reg_digest_next[21];   // sha_top.v(409)
    assign n3222 = rst ? 1'b0 : sha_reg_digest_next[20];   // sha_top.v(409)
    assign n3223 = rst ? 1'b0 : sha_reg_digest_next[19];   // sha_top.v(409)
    assign n3224 = rst ? 1'b0 : sha_reg_digest_next[18];   // sha_top.v(409)
    assign n3225 = rst ? 1'b0 : sha_reg_digest_next[17];   // sha_top.v(409)
    assign n3226 = rst ? 1'b0 : sha_reg_digest_next[16];   // sha_top.v(409)
    assign n3227 = rst ? 1'b0 : sha_reg_digest_next[15];   // sha_top.v(409)
    assign n3228 = rst ? 1'b0 : sha_reg_digest_next[14];   // sha_top.v(409)
    assign n3229 = rst ? 1'b0 : sha_reg_digest_next[13];   // sha_top.v(409)
    assign n3230 = rst ? 1'b0 : sha_reg_digest_next[12];   // sha_top.v(409)
    assign n3231 = rst ? 1'b0 : sha_reg_digest_next[11];   // sha_top.v(409)
    assign n3232 = rst ? 1'b0 : sha_reg_digest_next[10];   // sha_top.v(409)
    assign n3233 = rst ? 1'b0 : sha_reg_digest_next[9];   // sha_top.v(409)
    assign n3234 = rst ? 1'b0 : sha_reg_digest_next[8];   // sha_top.v(409)
    assign n3235 = rst ? 1'b0 : sha_reg_digest_next[7];   // sha_top.v(409)
    assign n3236 = rst ? 1'b0 : sha_reg_digest_next[6];   // sha_top.v(409)
    assign n3237 = rst ? 1'b0 : sha_reg_digest_next[5];   // sha_top.v(409)
    assign n3238 = rst ? 1'b0 : sha_reg_digest_next[4];   // sha_top.v(409)
    assign n3239 = rst ? 1'b0 : sha_reg_digest_next[3];   // sha_top.v(409)
    assign n3240 = rst ? 1'b0 : sha_reg_digest_next[2];   // sha_top.v(409)
    assign n3241 = rst ? 1'b0 : sha_reg_digest_next[1];   // sha_top.v(409)
    assign n3242 = rst ? 1'b0 : sha_reg_digest_next[0];   // sha_top.v(409)
    assign n3243 = rst ? 1'b0 : sha_core_ready;   // sha_top.v(409)
    VERIFIC_DFFRS i3165 (.d(n2531), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_state[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3166 (.d(n2532), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_state[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3167 (.d(n2533), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[5]));   // sha_top.v(410)
    VERIFIC_DFFRS i3168 (.d(n2534), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[4]));   // sha_top.v(410)
    VERIFIC_DFFRS i3169 (.d(n2535), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[3]));   // sha_top.v(410)
    VERIFIC_DFFRS i3170 (.d(n2536), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[2]));   // sha_top.v(410)
    VERIFIC_DFFRS i3171 (.d(n2537), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3172 (.d(n2538), .clk(clk), .s(1'b0), .r(1'b0), .q(byte_counter[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3173 (.d(n2539), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[511]));   // sha_top.v(410)
    VERIFIC_DFFRS i3174 (.d(n2540), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[510]));   // sha_top.v(410)
    VERIFIC_DFFRS i3175 (.d(n2541), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[509]));   // sha_top.v(410)
    VERIFIC_DFFRS i3176 (.d(n2542), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[508]));   // sha_top.v(410)
    VERIFIC_DFFRS i3177 (.d(n2543), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[507]));   // sha_top.v(410)
    VERIFIC_DFFRS i3178 (.d(n2544), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[506]));   // sha_top.v(410)
    VERIFIC_DFFRS i3179 (.d(n2545), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[505]));   // sha_top.v(410)
    VERIFIC_DFFRS i3180 (.d(n2546), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[504]));   // sha_top.v(410)
    VERIFIC_DFFRS i3181 (.d(n2547), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[503]));   // sha_top.v(410)
    VERIFIC_DFFRS i3182 (.d(n2548), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[502]));   // sha_top.v(410)
    VERIFIC_DFFRS i3183 (.d(n2549), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[501]));   // sha_top.v(410)
    VERIFIC_DFFRS i3184 (.d(n2550), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[500]));   // sha_top.v(410)
    VERIFIC_DFFRS i3185 (.d(n2551), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[499]));   // sha_top.v(410)
    VERIFIC_DFFRS i3186 (.d(n2552), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[498]));   // sha_top.v(410)
    VERIFIC_DFFRS i3187 (.d(n2553), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[497]));   // sha_top.v(410)
    VERIFIC_DFFRS i3188 (.d(n2554), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[496]));   // sha_top.v(410)
    VERIFIC_DFFRS i3189 (.d(n2555), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[495]));   // sha_top.v(410)
    VERIFIC_DFFRS i3190 (.d(n2556), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[494]));   // sha_top.v(410)
    VERIFIC_DFFRS i3191 (.d(n2557), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[493]));   // sha_top.v(410)
    VERIFIC_DFFRS i3192 (.d(n2558), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[492]));   // sha_top.v(410)
    VERIFIC_DFFRS i3193 (.d(n2559), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[491]));   // sha_top.v(410)
    VERIFIC_DFFRS i3194 (.d(n2560), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[490]));   // sha_top.v(410)
    VERIFIC_DFFRS i3195 (.d(n2561), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[489]));   // sha_top.v(410)
    VERIFIC_DFFRS i3196 (.d(n2562), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[488]));   // sha_top.v(410)
    VERIFIC_DFFRS i3197 (.d(n2563), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[487]));   // sha_top.v(410)
    VERIFIC_DFFRS i3198 (.d(n2564), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[486]));   // sha_top.v(410)
    VERIFIC_DFFRS i3199 (.d(n2565), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[485]));   // sha_top.v(410)
    VERIFIC_DFFRS i3200 (.d(n2566), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[484]));   // sha_top.v(410)
    VERIFIC_DFFRS i3201 (.d(n2567), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[483]));   // sha_top.v(410)
    VERIFIC_DFFRS i3202 (.d(n2568), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[482]));   // sha_top.v(410)
    VERIFIC_DFFRS i3203 (.d(n2569), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[481]));   // sha_top.v(410)
    VERIFIC_DFFRS i3204 (.d(n2570), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[480]));   // sha_top.v(410)
    VERIFIC_DFFRS i3205 (.d(n2571), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[479]));   // sha_top.v(410)
    VERIFIC_DFFRS i3206 (.d(n2572), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[478]));   // sha_top.v(410)
    VERIFIC_DFFRS i3207 (.d(n2573), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[477]));   // sha_top.v(410)
    VERIFIC_DFFRS i3208 (.d(n2574), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[476]));   // sha_top.v(410)
    VERIFIC_DFFRS i3209 (.d(n2575), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[475]));   // sha_top.v(410)
    VERIFIC_DFFRS i3210 (.d(n2576), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[474]));   // sha_top.v(410)
    VERIFIC_DFFRS i3211 (.d(n2577), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[473]));   // sha_top.v(410)
    VERIFIC_DFFRS i3212 (.d(n2578), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[472]));   // sha_top.v(410)
    VERIFIC_DFFRS i3213 (.d(n2579), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[471]));   // sha_top.v(410)
    VERIFIC_DFFRS i3214 (.d(n2580), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[470]));   // sha_top.v(410)
    VERIFIC_DFFRS i3215 (.d(n2581), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[469]));   // sha_top.v(410)
    VERIFIC_DFFRS i3216 (.d(n2582), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[468]));   // sha_top.v(410)
    VERIFIC_DFFRS i3217 (.d(n2583), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[467]));   // sha_top.v(410)
    VERIFIC_DFFRS i3218 (.d(n2584), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[466]));   // sha_top.v(410)
    VERIFIC_DFFRS i3219 (.d(n2585), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[465]));   // sha_top.v(410)
    VERIFIC_DFFRS i3220 (.d(n2586), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[464]));   // sha_top.v(410)
    VERIFIC_DFFRS i3221 (.d(n2587), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[463]));   // sha_top.v(410)
    VERIFIC_DFFRS i3222 (.d(n2588), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[462]));   // sha_top.v(410)
    VERIFIC_DFFRS i3223 (.d(n2589), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[461]));   // sha_top.v(410)
    VERIFIC_DFFRS i3224 (.d(n2590), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[460]));   // sha_top.v(410)
    VERIFIC_DFFRS i3225 (.d(n2591), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[459]));   // sha_top.v(410)
    VERIFIC_DFFRS i3226 (.d(n2592), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[458]));   // sha_top.v(410)
    VERIFIC_DFFRS i3227 (.d(n2593), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[457]));   // sha_top.v(410)
    VERIFIC_DFFRS i3228 (.d(n2594), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[456]));   // sha_top.v(410)
    VERIFIC_DFFRS i3229 (.d(n2595), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[455]));   // sha_top.v(410)
    VERIFIC_DFFRS i3230 (.d(n2596), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[454]));   // sha_top.v(410)
    VERIFIC_DFFRS i3231 (.d(n2597), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[453]));   // sha_top.v(410)
    VERIFIC_DFFRS i3232 (.d(n2598), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[452]));   // sha_top.v(410)
    VERIFIC_DFFRS i3233 (.d(n2599), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[451]));   // sha_top.v(410)
    VERIFIC_DFFRS i3234 (.d(n2600), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[450]));   // sha_top.v(410)
    VERIFIC_DFFRS i3235 (.d(n2601), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[449]));   // sha_top.v(410)
    VERIFIC_DFFRS i3236 (.d(n2602), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[448]));   // sha_top.v(410)
    VERIFIC_DFFRS i3237 (.d(n2603), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[447]));   // sha_top.v(410)
    VERIFIC_DFFRS i3238 (.d(n2604), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[446]));   // sha_top.v(410)
    VERIFIC_DFFRS i3239 (.d(n2605), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[445]));   // sha_top.v(410)
    VERIFIC_DFFRS i3240 (.d(n2606), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[444]));   // sha_top.v(410)
    VERIFIC_DFFRS i3241 (.d(n2607), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[443]));   // sha_top.v(410)
    VERIFIC_DFFRS i3242 (.d(n2608), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[442]));   // sha_top.v(410)
    VERIFIC_DFFRS i3243 (.d(n2609), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[441]));   // sha_top.v(410)
    VERIFIC_DFFRS i3244 (.d(n2610), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[440]));   // sha_top.v(410)
    VERIFIC_DFFRS i3245 (.d(n2611), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[439]));   // sha_top.v(410)
    VERIFIC_DFFRS i3246 (.d(n2612), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[438]));   // sha_top.v(410)
    VERIFIC_DFFRS i3247 (.d(n2613), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[437]));   // sha_top.v(410)
    VERIFIC_DFFRS i3248 (.d(n2614), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[436]));   // sha_top.v(410)
    VERIFIC_DFFRS i3249 (.d(n2615), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[435]));   // sha_top.v(410)
    VERIFIC_DFFRS i3250 (.d(n2616), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[434]));   // sha_top.v(410)
    VERIFIC_DFFRS i3251 (.d(n2617), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[433]));   // sha_top.v(410)
    VERIFIC_DFFRS i3252 (.d(n2618), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[432]));   // sha_top.v(410)
    VERIFIC_DFFRS i3253 (.d(n2619), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[431]));   // sha_top.v(410)
    VERIFIC_DFFRS i3254 (.d(n2620), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[430]));   // sha_top.v(410)
    VERIFIC_DFFRS i3255 (.d(n2621), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[429]));   // sha_top.v(410)
    VERIFIC_DFFRS i3256 (.d(n2622), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[428]));   // sha_top.v(410)
    VERIFIC_DFFRS i3257 (.d(n2623), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[427]));   // sha_top.v(410)
    VERIFIC_DFFRS i3258 (.d(n2624), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[426]));   // sha_top.v(410)
    VERIFIC_DFFRS i3259 (.d(n2625), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[425]));   // sha_top.v(410)
    VERIFIC_DFFRS i3260 (.d(n2626), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[424]));   // sha_top.v(410)
    VERIFIC_DFFRS i3261 (.d(n2627), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[423]));   // sha_top.v(410)
    VERIFIC_DFFRS i3262 (.d(n2628), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[422]));   // sha_top.v(410)
    VERIFIC_DFFRS i3263 (.d(n2629), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[421]));   // sha_top.v(410)
    VERIFIC_DFFRS i3264 (.d(n2630), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[420]));   // sha_top.v(410)
    VERIFIC_DFFRS i3265 (.d(n2631), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[419]));   // sha_top.v(410)
    VERIFIC_DFFRS i3266 (.d(n2632), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[418]));   // sha_top.v(410)
    VERIFIC_DFFRS i3267 (.d(n2633), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[417]));   // sha_top.v(410)
    VERIFIC_DFFRS i3268 (.d(n2634), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[416]));   // sha_top.v(410)
    VERIFIC_DFFRS i3269 (.d(n2635), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[415]));   // sha_top.v(410)
    VERIFIC_DFFRS i3270 (.d(n2636), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[414]));   // sha_top.v(410)
    VERIFIC_DFFRS i3271 (.d(n2637), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[413]));   // sha_top.v(410)
    VERIFIC_DFFRS i3272 (.d(n2638), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[412]));   // sha_top.v(410)
    VERIFIC_DFFRS i3273 (.d(n2639), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[411]));   // sha_top.v(410)
    VERIFIC_DFFRS i3274 (.d(n2640), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[410]));   // sha_top.v(410)
    VERIFIC_DFFRS i3275 (.d(n2641), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[409]));   // sha_top.v(410)
    VERIFIC_DFFRS i3276 (.d(n2642), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[408]));   // sha_top.v(410)
    VERIFIC_DFFRS i3277 (.d(n2643), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[407]));   // sha_top.v(410)
    VERIFIC_DFFRS i3278 (.d(n2644), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[406]));   // sha_top.v(410)
    VERIFIC_DFFRS i3279 (.d(n2645), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[405]));   // sha_top.v(410)
    VERIFIC_DFFRS i3280 (.d(n2646), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[404]));   // sha_top.v(410)
    VERIFIC_DFFRS i3281 (.d(n2647), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[403]));   // sha_top.v(410)
    VERIFIC_DFFRS i3282 (.d(n2648), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[402]));   // sha_top.v(410)
    VERIFIC_DFFRS i3283 (.d(n2649), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[401]));   // sha_top.v(410)
    VERIFIC_DFFRS i3284 (.d(n2650), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[400]));   // sha_top.v(410)
    VERIFIC_DFFRS i3285 (.d(n2651), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[399]));   // sha_top.v(410)
    VERIFIC_DFFRS i3286 (.d(n2652), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[398]));   // sha_top.v(410)
    VERIFIC_DFFRS i3287 (.d(n2653), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[397]));   // sha_top.v(410)
    VERIFIC_DFFRS i3288 (.d(n2654), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[396]));   // sha_top.v(410)
    VERIFIC_DFFRS i3289 (.d(n2655), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[395]));   // sha_top.v(410)
    VERIFIC_DFFRS i3290 (.d(n2656), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[394]));   // sha_top.v(410)
    VERIFIC_DFFRS i3291 (.d(n2657), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[393]));   // sha_top.v(410)
    VERIFIC_DFFRS i3292 (.d(n2658), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[392]));   // sha_top.v(410)
    VERIFIC_DFFRS i3293 (.d(n2659), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[391]));   // sha_top.v(410)
    VERIFIC_DFFRS i3294 (.d(n2660), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[390]));   // sha_top.v(410)
    VERIFIC_DFFRS i3295 (.d(n2661), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[389]));   // sha_top.v(410)
    VERIFIC_DFFRS i3296 (.d(n2662), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[388]));   // sha_top.v(410)
    VERIFIC_DFFRS i3297 (.d(n2663), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[387]));   // sha_top.v(410)
    VERIFIC_DFFRS i3298 (.d(n2664), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[386]));   // sha_top.v(410)
    VERIFIC_DFFRS i3299 (.d(n2665), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[385]));   // sha_top.v(410)
    VERIFIC_DFFRS i3300 (.d(n2666), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[384]));   // sha_top.v(410)
    VERIFIC_DFFRS i3301 (.d(n2667), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[383]));   // sha_top.v(410)
    VERIFIC_DFFRS i3302 (.d(n2668), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[382]));   // sha_top.v(410)
    VERIFIC_DFFRS i3303 (.d(n2669), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[381]));   // sha_top.v(410)
    VERIFIC_DFFRS i3304 (.d(n2670), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[380]));   // sha_top.v(410)
    VERIFIC_DFFRS i3305 (.d(n2671), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[379]));   // sha_top.v(410)
    VERIFIC_DFFRS i3306 (.d(n2672), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[378]));   // sha_top.v(410)
    VERIFIC_DFFRS i3307 (.d(n2673), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[377]));   // sha_top.v(410)
    VERIFIC_DFFRS i3308 (.d(n2674), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[376]));   // sha_top.v(410)
    VERIFIC_DFFRS i3309 (.d(n2675), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[375]));   // sha_top.v(410)
    VERIFIC_DFFRS i3310 (.d(n2676), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[374]));   // sha_top.v(410)
    VERIFIC_DFFRS i3311 (.d(n2677), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[373]));   // sha_top.v(410)
    VERIFIC_DFFRS i3312 (.d(n2678), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[372]));   // sha_top.v(410)
    VERIFIC_DFFRS i3313 (.d(n2679), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[371]));   // sha_top.v(410)
    VERIFIC_DFFRS i3314 (.d(n2680), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[370]));   // sha_top.v(410)
    VERIFIC_DFFRS i3315 (.d(n2681), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[369]));   // sha_top.v(410)
    VERIFIC_DFFRS i3316 (.d(n2682), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[368]));   // sha_top.v(410)
    VERIFIC_DFFRS i3317 (.d(n2683), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[367]));   // sha_top.v(410)
    VERIFIC_DFFRS i3318 (.d(n2684), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[366]));   // sha_top.v(410)
    VERIFIC_DFFRS i3319 (.d(n2685), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[365]));   // sha_top.v(410)
    VERIFIC_DFFRS i3320 (.d(n2686), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[364]));   // sha_top.v(410)
    VERIFIC_DFFRS i3321 (.d(n2687), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[363]));   // sha_top.v(410)
    VERIFIC_DFFRS i3322 (.d(n2688), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[362]));   // sha_top.v(410)
    VERIFIC_DFFRS i3323 (.d(n2689), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[361]));   // sha_top.v(410)
    VERIFIC_DFFRS i3324 (.d(n2690), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[360]));   // sha_top.v(410)
    VERIFIC_DFFRS i3325 (.d(n2691), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[359]));   // sha_top.v(410)
    VERIFIC_DFFRS i3326 (.d(n2692), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[358]));   // sha_top.v(410)
    VERIFIC_DFFRS i3327 (.d(n2693), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[357]));   // sha_top.v(410)
    VERIFIC_DFFRS i3328 (.d(n2694), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[356]));   // sha_top.v(410)
    VERIFIC_DFFRS i3329 (.d(n2695), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[355]));   // sha_top.v(410)
    VERIFIC_DFFRS i3330 (.d(n2696), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[354]));   // sha_top.v(410)
    VERIFIC_DFFRS i3331 (.d(n2697), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[353]));   // sha_top.v(410)
    VERIFIC_DFFRS i3332 (.d(n2698), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[352]));   // sha_top.v(410)
    VERIFIC_DFFRS i3333 (.d(n2699), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[351]));   // sha_top.v(410)
    VERIFIC_DFFRS i3334 (.d(n2700), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[350]));   // sha_top.v(410)
    VERIFIC_DFFRS i3335 (.d(n2701), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[349]));   // sha_top.v(410)
    VERIFIC_DFFRS i3336 (.d(n2702), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[348]));   // sha_top.v(410)
    VERIFIC_DFFRS i3337 (.d(n2703), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[347]));   // sha_top.v(410)
    VERIFIC_DFFRS i3338 (.d(n2704), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[346]));   // sha_top.v(410)
    VERIFIC_DFFRS i3339 (.d(n2705), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[345]));   // sha_top.v(410)
    VERIFIC_DFFRS i3340 (.d(n2706), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[344]));   // sha_top.v(410)
    VERIFIC_DFFRS i3341 (.d(n2707), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[343]));   // sha_top.v(410)
    VERIFIC_DFFRS i3342 (.d(n2708), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[342]));   // sha_top.v(410)
    VERIFIC_DFFRS i3343 (.d(n2709), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[341]));   // sha_top.v(410)
    VERIFIC_DFFRS i3344 (.d(n2710), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[340]));   // sha_top.v(410)
    VERIFIC_DFFRS i3345 (.d(n2711), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[339]));   // sha_top.v(410)
    VERIFIC_DFFRS i3346 (.d(n2712), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[338]));   // sha_top.v(410)
    VERIFIC_DFFRS i3347 (.d(n2713), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[337]));   // sha_top.v(410)
    VERIFIC_DFFRS i3348 (.d(n2714), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[336]));   // sha_top.v(410)
    VERIFIC_DFFRS i3349 (.d(n2715), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[335]));   // sha_top.v(410)
    VERIFIC_DFFRS i3350 (.d(n2716), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[334]));   // sha_top.v(410)
    VERIFIC_DFFRS i3351 (.d(n2717), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[333]));   // sha_top.v(410)
    VERIFIC_DFFRS i3352 (.d(n2718), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[332]));   // sha_top.v(410)
    VERIFIC_DFFRS i3353 (.d(n2719), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[331]));   // sha_top.v(410)
    VERIFIC_DFFRS i3354 (.d(n2720), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[330]));   // sha_top.v(410)
    VERIFIC_DFFRS i3355 (.d(n2721), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[329]));   // sha_top.v(410)
    VERIFIC_DFFRS i3356 (.d(n2722), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[328]));   // sha_top.v(410)
    VERIFIC_DFFRS i3357 (.d(n2723), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[327]));   // sha_top.v(410)
    VERIFIC_DFFRS i3358 (.d(n2724), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[326]));   // sha_top.v(410)
    VERIFIC_DFFRS i3359 (.d(n2725), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[325]));   // sha_top.v(410)
    VERIFIC_DFFRS i3360 (.d(n2726), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[324]));   // sha_top.v(410)
    VERIFIC_DFFRS i3361 (.d(n2727), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[323]));   // sha_top.v(410)
    VERIFIC_DFFRS i3362 (.d(n2728), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[322]));   // sha_top.v(410)
    VERIFIC_DFFRS i3363 (.d(n2729), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[321]));   // sha_top.v(410)
    VERIFIC_DFFRS i3364 (.d(n2730), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[320]));   // sha_top.v(410)
    VERIFIC_DFFRS i3365 (.d(n2731), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[319]));   // sha_top.v(410)
    VERIFIC_DFFRS i3366 (.d(n2732), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[318]));   // sha_top.v(410)
    VERIFIC_DFFRS i3367 (.d(n2733), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[317]));   // sha_top.v(410)
    VERIFIC_DFFRS i3368 (.d(n2734), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[316]));   // sha_top.v(410)
    VERIFIC_DFFRS i3369 (.d(n2735), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[315]));   // sha_top.v(410)
    VERIFIC_DFFRS i3370 (.d(n2736), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[314]));   // sha_top.v(410)
    VERIFIC_DFFRS i3371 (.d(n2737), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[313]));   // sha_top.v(410)
    VERIFIC_DFFRS i3372 (.d(n2738), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[312]));   // sha_top.v(410)
    VERIFIC_DFFRS i3373 (.d(n2739), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[311]));   // sha_top.v(410)
    VERIFIC_DFFRS i3374 (.d(n2740), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[310]));   // sha_top.v(410)
    VERIFIC_DFFRS i3375 (.d(n2741), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[309]));   // sha_top.v(410)
    VERIFIC_DFFRS i3376 (.d(n2742), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[308]));   // sha_top.v(410)
    VERIFIC_DFFRS i3377 (.d(n2743), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[307]));   // sha_top.v(410)
    VERIFIC_DFFRS i3378 (.d(n2744), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[306]));   // sha_top.v(410)
    VERIFIC_DFFRS i3379 (.d(n2745), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[305]));   // sha_top.v(410)
    VERIFIC_DFFRS i3380 (.d(n2746), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[304]));   // sha_top.v(410)
    VERIFIC_DFFRS i3381 (.d(n2747), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[303]));   // sha_top.v(410)
    VERIFIC_DFFRS i3382 (.d(n2748), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[302]));   // sha_top.v(410)
    VERIFIC_DFFRS i3383 (.d(n2749), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[301]));   // sha_top.v(410)
    VERIFIC_DFFRS i3384 (.d(n2750), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[300]));   // sha_top.v(410)
    VERIFIC_DFFRS i3385 (.d(n2751), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[299]));   // sha_top.v(410)
    VERIFIC_DFFRS i3386 (.d(n2752), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[298]));   // sha_top.v(410)
    VERIFIC_DFFRS i3387 (.d(n2753), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[297]));   // sha_top.v(410)
    VERIFIC_DFFRS i3388 (.d(n2754), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[296]));   // sha_top.v(410)
    VERIFIC_DFFRS i3389 (.d(n2755), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[295]));   // sha_top.v(410)
    VERIFIC_DFFRS i3390 (.d(n2756), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[294]));   // sha_top.v(410)
    VERIFIC_DFFRS i3391 (.d(n2757), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[293]));   // sha_top.v(410)
    VERIFIC_DFFRS i3392 (.d(n2758), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[292]));   // sha_top.v(410)
    VERIFIC_DFFRS i3393 (.d(n2759), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[291]));   // sha_top.v(410)
    VERIFIC_DFFRS i3394 (.d(n2760), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[290]));   // sha_top.v(410)
    VERIFIC_DFFRS i3395 (.d(n2761), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[289]));   // sha_top.v(410)
    VERIFIC_DFFRS i3396 (.d(n2762), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[288]));   // sha_top.v(410)
    VERIFIC_DFFRS i3397 (.d(n2763), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[287]));   // sha_top.v(410)
    VERIFIC_DFFRS i3398 (.d(n2764), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[286]));   // sha_top.v(410)
    VERIFIC_DFFRS i3399 (.d(n2765), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[285]));   // sha_top.v(410)
    VERIFIC_DFFRS i3400 (.d(n2766), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[284]));   // sha_top.v(410)
    VERIFIC_DFFRS i3401 (.d(n2767), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[283]));   // sha_top.v(410)
    VERIFIC_DFFRS i3402 (.d(n2768), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[282]));   // sha_top.v(410)
    VERIFIC_DFFRS i3403 (.d(n2769), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[281]));   // sha_top.v(410)
    VERIFIC_DFFRS i3404 (.d(n2770), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[280]));   // sha_top.v(410)
    VERIFIC_DFFRS i3405 (.d(n2771), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[279]));   // sha_top.v(410)
    VERIFIC_DFFRS i3406 (.d(n2772), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[278]));   // sha_top.v(410)
    VERIFIC_DFFRS i3407 (.d(n2773), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[277]));   // sha_top.v(410)
    VERIFIC_DFFRS i3408 (.d(n2774), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[276]));   // sha_top.v(410)
    VERIFIC_DFFRS i3409 (.d(n2775), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[275]));   // sha_top.v(410)
    VERIFIC_DFFRS i3410 (.d(n2776), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[274]));   // sha_top.v(410)
    VERIFIC_DFFRS i3411 (.d(n2777), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[273]));   // sha_top.v(410)
    VERIFIC_DFFRS i3412 (.d(n2778), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[272]));   // sha_top.v(410)
    VERIFIC_DFFRS i3413 (.d(n2779), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[271]));   // sha_top.v(410)
    VERIFIC_DFFRS i3414 (.d(n2780), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[270]));   // sha_top.v(410)
    VERIFIC_DFFRS i3415 (.d(n2781), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[269]));   // sha_top.v(410)
    VERIFIC_DFFRS i3416 (.d(n2782), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[268]));   // sha_top.v(410)
    VERIFIC_DFFRS i3417 (.d(n2783), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[267]));   // sha_top.v(410)
    VERIFIC_DFFRS i3418 (.d(n2784), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[266]));   // sha_top.v(410)
    VERIFIC_DFFRS i3419 (.d(n2785), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[265]));   // sha_top.v(410)
    VERIFIC_DFFRS i3420 (.d(n2786), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[264]));   // sha_top.v(410)
    VERIFIC_DFFRS i3421 (.d(n2787), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[263]));   // sha_top.v(410)
    VERIFIC_DFFRS i3422 (.d(n2788), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[262]));   // sha_top.v(410)
    VERIFIC_DFFRS i3423 (.d(n2789), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[261]));   // sha_top.v(410)
    VERIFIC_DFFRS i3424 (.d(n2790), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[260]));   // sha_top.v(410)
    VERIFIC_DFFRS i3425 (.d(n2791), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[259]));   // sha_top.v(410)
    VERIFIC_DFFRS i3426 (.d(n2792), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[258]));   // sha_top.v(410)
    VERIFIC_DFFRS i3427 (.d(n2793), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[257]));   // sha_top.v(410)
    VERIFIC_DFFRS i3428 (.d(n2794), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[256]));   // sha_top.v(410)
    VERIFIC_DFFRS i3429 (.d(n2795), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[255]));   // sha_top.v(410)
    VERIFIC_DFFRS i3430 (.d(n2796), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[254]));   // sha_top.v(410)
    VERIFIC_DFFRS i3431 (.d(n2797), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[253]));   // sha_top.v(410)
    VERIFIC_DFFRS i3432 (.d(n2798), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[252]));   // sha_top.v(410)
    VERIFIC_DFFRS i3433 (.d(n2799), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[251]));   // sha_top.v(410)
    VERIFIC_DFFRS i3434 (.d(n2800), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[250]));   // sha_top.v(410)
    VERIFIC_DFFRS i3435 (.d(n2801), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[249]));   // sha_top.v(410)
    VERIFIC_DFFRS i3436 (.d(n2802), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[248]));   // sha_top.v(410)
    VERIFIC_DFFRS i3437 (.d(n2803), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[247]));   // sha_top.v(410)
    VERIFIC_DFFRS i3438 (.d(n2804), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[246]));   // sha_top.v(410)
    VERIFIC_DFFRS i3439 (.d(n2805), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[245]));   // sha_top.v(410)
    VERIFIC_DFFRS i3440 (.d(n2806), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[244]));   // sha_top.v(410)
    VERIFIC_DFFRS i3441 (.d(n2807), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[243]));   // sha_top.v(410)
    VERIFIC_DFFRS i3442 (.d(n2808), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[242]));   // sha_top.v(410)
    VERIFIC_DFFRS i3443 (.d(n2809), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[241]));   // sha_top.v(410)
    VERIFIC_DFFRS i3444 (.d(n2810), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[240]));   // sha_top.v(410)
    VERIFIC_DFFRS i3445 (.d(n2811), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[239]));   // sha_top.v(410)
    VERIFIC_DFFRS i3446 (.d(n2812), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[238]));   // sha_top.v(410)
    VERIFIC_DFFRS i3447 (.d(n2813), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[237]));   // sha_top.v(410)
    VERIFIC_DFFRS i3448 (.d(n2814), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[236]));   // sha_top.v(410)
    VERIFIC_DFFRS i3449 (.d(n2815), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[235]));   // sha_top.v(410)
    VERIFIC_DFFRS i3450 (.d(n2816), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[234]));   // sha_top.v(410)
    VERIFIC_DFFRS i3451 (.d(n2817), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[233]));   // sha_top.v(410)
    VERIFIC_DFFRS i3452 (.d(n2818), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[232]));   // sha_top.v(410)
    VERIFIC_DFFRS i3453 (.d(n2819), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[231]));   // sha_top.v(410)
    VERIFIC_DFFRS i3454 (.d(n2820), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[230]));   // sha_top.v(410)
    VERIFIC_DFFRS i3455 (.d(n2821), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[229]));   // sha_top.v(410)
    VERIFIC_DFFRS i3456 (.d(n2822), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[228]));   // sha_top.v(410)
    VERIFIC_DFFRS i3457 (.d(n2823), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[227]));   // sha_top.v(410)
    VERIFIC_DFFRS i3458 (.d(n2824), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[226]));   // sha_top.v(410)
    VERIFIC_DFFRS i3459 (.d(n2825), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[225]));   // sha_top.v(410)
    VERIFIC_DFFRS i3460 (.d(n2826), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[224]));   // sha_top.v(410)
    VERIFIC_DFFRS i3461 (.d(n2827), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[223]));   // sha_top.v(410)
    VERIFIC_DFFRS i3462 (.d(n2828), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[222]));   // sha_top.v(410)
    VERIFIC_DFFRS i3463 (.d(n2829), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[221]));   // sha_top.v(410)
    VERIFIC_DFFRS i3464 (.d(n2830), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[220]));   // sha_top.v(410)
    VERIFIC_DFFRS i3465 (.d(n2831), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[219]));   // sha_top.v(410)
    VERIFIC_DFFRS i3466 (.d(n2832), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[218]));   // sha_top.v(410)
    VERIFIC_DFFRS i3467 (.d(n2833), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[217]));   // sha_top.v(410)
    VERIFIC_DFFRS i3468 (.d(n2834), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[216]));   // sha_top.v(410)
    VERIFIC_DFFRS i3469 (.d(n2835), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[215]));   // sha_top.v(410)
    VERIFIC_DFFRS i3470 (.d(n2836), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[214]));   // sha_top.v(410)
    VERIFIC_DFFRS i3471 (.d(n2837), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[213]));   // sha_top.v(410)
    VERIFIC_DFFRS i3472 (.d(n2838), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[212]));   // sha_top.v(410)
    VERIFIC_DFFRS i3473 (.d(n2839), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[211]));   // sha_top.v(410)
    VERIFIC_DFFRS i3474 (.d(n2840), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[210]));   // sha_top.v(410)
    VERIFIC_DFFRS i3475 (.d(n2841), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[209]));   // sha_top.v(410)
    VERIFIC_DFFRS i3476 (.d(n2842), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[208]));   // sha_top.v(410)
    VERIFIC_DFFRS i3477 (.d(n2843), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[207]));   // sha_top.v(410)
    VERIFIC_DFFRS i3478 (.d(n2844), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[206]));   // sha_top.v(410)
    VERIFIC_DFFRS i3479 (.d(n2845), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[205]));   // sha_top.v(410)
    VERIFIC_DFFRS i3480 (.d(n2846), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[204]));   // sha_top.v(410)
    VERIFIC_DFFRS i3481 (.d(n2847), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[203]));   // sha_top.v(410)
    VERIFIC_DFFRS i3482 (.d(n2848), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[202]));   // sha_top.v(410)
    VERIFIC_DFFRS i3483 (.d(n2849), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[201]));   // sha_top.v(410)
    VERIFIC_DFFRS i3484 (.d(n2850), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[200]));   // sha_top.v(410)
    VERIFIC_DFFRS i3485 (.d(n2851), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[199]));   // sha_top.v(410)
    VERIFIC_DFFRS i3486 (.d(n2852), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[198]));   // sha_top.v(410)
    VERIFIC_DFFRS i3487 (.d(n2853), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[197]));   // sha_top.v(410)
    VERIFIC_DFFRS i3488 (.d(n2854), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[196]));   // sha_top.v(410)
    VERIFIC_DFFRS i3489 (.d(n2855), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[195]));   // sha_top.v(410)
    VERIFIC_DFFRS i3490 (.d(n2856), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[194]));   // sha_top.v(410)
    VERIFIC_DFFRS i3491 (.d(n2857), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[193]));   // sha_top.v(410)
    VERIFIC_DFFRS i3492 (.d(n2858), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[192]));   // sha_top.v(410)
    VERIFIC_DFFRS i3493 (.d(n2859), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[191]));   // sha_top.v(410)
    VERIFIC_DFFRS i3494 (.d(n2860), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[190]));   // sha_top.v(410)
    VERIFIC_DFFRS i3495 (.d(n2861), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[189]));   // sha_top.v(410)
    VERIFIC_DFFRS i3496 (.d(n2862), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[188]));   // sha_top.v(410)
    VERIFIC_DFFRS i3497 (.d(n2863), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[187]));   // sha_top.v(410)
    VERIFIC_DFFRS i3498 (.d(n2864), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[186]));   // sha_top.v(410)
    VERIFIC_DFFRS i3499 (.d(n2865), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[185]));   // sha_top.v(410)
    VERIFIC_DFFRS i3500 (.d(n2866), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[184]));   // sha_top.v(410)
    VERIFIC_DFFRS i3501 (.d(n2867), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[183]));   // sha_top.v(410)
    VERIFIC_DFFRS i3502 (.d(n2868), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[182]));   // sha_top.v(410)
    VERIFIC_DFFRS i3503 (.d(n2869), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[181]));   // sha_top.v(410)
    VERIFIC_DFFRS i3504 (.d(n2870), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[180]));   // sha_top.v(410)
    VERIFIC_DFFRS i3505 (.d(n2871), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[179]));   // sha_top.v(410)
    VERIFIC_DFFRS i3506 (.d(n2872), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[178]));   // sha_top.v(410)
    VERIFIC_DFFRS i3507 (.d(n2873), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[177]));   // sha_top.v(410)
    VERIFIC_DFFRS i3508 (.d(n2874), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[176]));   // sha_top.v(410)
    VERIFIC_DFFRS i3509 (.d(n2875), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[175]));   // sha_top.v(410)
    VERIFIC_DFFRS i3510 (.d(n2876), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[174]));   // sha_top.v(410)
    VERIFIC_DFFRS i3511 (.d(n2877), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[173]));   // sha_top.v(410)
    VERIFIC_DFFRS i3512 (.d(n2878), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[172]));   // sha_top.v(410)
    VERIFIC_DFFRS i3513 (.d(n2879), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[171]));   // sha_top.v(410)
    VERIFIC_DFFRS i3514 (.d(n2880), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[170]));   // sha_top.v(410)
    VERIFIC_DFFRS i3515 (.d(n2881), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[169]));   // sha_top.v(410)
    VERIFIC_DFFRS i3516 (.d(n2882), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[168]));   // sha_top.v(410)
    VERIFIC_DFFRS i3517 (.d(n2883), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[167]));   // sha_top.v(410)
    VERIFIC_DFFRS i3518 (.d(n2884), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[166]));   // sha_top.v(410)
    VERIFIC_DFFRS i3519 (.d(n2885), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[165]));   // sha_top.v(410)
    VERIFIC_DFFRS i3520 (.d(n2886), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[164]));   // sha_top.v(410)
    VERIFIC_DFFRS i3521 (.d(n2887), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[163]));   // sha_top.v(410)
    VERIFIC_DFFRS i3522 (.d(n2888), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[162]));   // sha_top.v(410)
    VERIFIC_DFFRS i3523 (.d(n2889), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[161]));   // sha_top.v(410)
    VERIFIC_DFFRS i3524 (.d(n2890), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[160]));   // sha_top.v(410)
    VERIFIC_DFFRS i3525 (.d(n2891), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[159]));   // sha_top.v(410)
    VERIFIC_DFFRS i3526 (.d(n2892), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[158]));   // sha_top.v(410)
    VERIFIC_DFFRS i3527 (.d(n2893), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[157]));   // sha_top.v(410)
    VERIFIC_DFFRS i3528 (.d(n2894), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[156]));   // sha_top.v(410)
    VERIFIC_DFFRS i3529 (.d(n2895), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[155]));   // sha_top.v(410)
    VERIFIC_DFFRS i3530 (.d(n2896), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[154]));   // sha_top.v(410)
    VERIFIC_DFFRS i3531 (.d(n2897), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[153]));   // sha_top.v(410)
    VERIFIC_DFFRS i3532 (.d(n2898), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[152]));   // sha_top.v(410)
    VERIFIC_DFFRS i3533 (.d(n2899), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[151]));   // sha_top.v(410)
    VERIFIC_DFFRS i3534 (.d(n2900), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[150]));   // sha_top.v(410)
    VERIFIC_DFFRS i3535 (.d(n2901), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[149]));   // sha_top.v(410)
    VERIFIC_DFFRS i3536 (.d(n2902), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[148]));   // sha_top.v(410)
    VERIFIC_DFFRS i3537 (.d(n2903), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[147]));   // sha_top.v(410)
    VERIFIC_DFFRS i3538 (.d(n2904), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[146]));   // sha_top.v(410)
    VERIFIC_DFFRS i3539 (.d(n2905), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[145]));   // sha_top.v(410)
    VERIFIC_DFFRS i3540 (.d(n2906), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[144]));   // sha_top.v(410)
    VERIFIC_DFFRS i3541 (.d(n2907), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[143]));   // sha_top.v(410)
    VERIFIC_DFFRS i3542 (.d(n2908), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[142]));   // sha_top.v(410)
    VERIFIC_DFFRS i3543 (.d(n2909), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[141]));   // sha_top.v(410)
    VERIFIC_DFFRS i3544 (.d(n2910), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[140]));   // sha_top.v(410)
    VERIFIC_DFFRS i3545 (.d(n2911), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[139]));   // sha_top.v(410)
    VERIFIC_DFFRS i3546 (.d(n2912), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[138]));   // sha_top.v(410)
    VERIFIC_DFFRS i3547 (.d(n2913), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[137]));   // sha_top.v(410)
    VERIFIC_DFFRS i3548 (.d(n2914), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[136]));   // sha_top.v(410)
    VERIFIC_DFFRS i3549 (.d(n2915), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[135]));   // sha_top.v(410)
    VERIFIC_DFFRS i3550 (.d(n2916), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[134]));   // sha_top.v(410)
    VERIFIC_DFFRS i3551 (.d(n2917), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[133]));   // sha_top.v(410)
    VERIFIC_DFFRS i3552 (.d(n2918), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[132]));   // sha_top.v(410)
    VERIFIC_DFFRS i3553 (.d(n2919), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[131]));   // sha_top.v(410)
    VERIFIC_DFFRS i3554 (.d(n2920), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[130]));   // sha_top.v(410)
    VERIFIC_DFFRS i3555 (.d(n2921), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[129]));   // sha_top.v(410)
    VERIFIC_DFFRS i3556 (.d(n2922), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[128]));   // sha_top.v(410)
    VERIFIC_DFFRS i3557 (.d(n2923), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[127]));   // sha_top.v(410)
    VERIFIC_DFFRS i3558 (.d(n2924), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[126]));   // sha_top.v(410)
    VERIFIC_DFFRS i3559 (.d(n2925), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[125]));   // sha_top.v(410)
    VERIFIC_DFFRS i3560 (.d(n2926), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[124]));   // sha_top.v(410)
    VERIFIC_DFFRS i3561 (.d(n2927), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[123]));   // sha_top.v(410)
    VERIFIC_DFFRS i3562 (.d(n2928), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[122]));   // sha_top.v(410)
    VERIFIC_DFFRS i3563 (.d(n2929), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[121]));   // sha_top.v(410)
    VERIFIC_DFFRS i3564 (.d(n2930), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[120]));   // sha_top.v(410)
    VERIFIC_DFFRS i3565 (.d(n2931), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[119]));   // sha_top.v(410)
    VERIFIC_DFFRS i3566 (.d(n2932), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[118]));   // sha_top.v(410)
    VERIFIC_DFFRS i3567 (.d(n2933), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[117]));   // sha_top.v(410)
    VERIFIC_DFFRS i3568 (.d(n2934), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[116]));   // sha_top.v(410)
    VERIFIC_DFFRS i3569 (.d(n2935), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[115]));   // sha_top.v(410)
    VERIFIC_DFFRS i3570 (.d(n2936), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[114]));   // sha_top.v(410)
    VERIFIC_DFFRS i3571 (.d(n2937), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[113]));   // sha_top.v(410)
    VERIFIC_DFFRS i3572 (.d(n2938), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[112]));   // sha_top.v(410)
    VERIFIC_DFFRS i3573 (.d(n2939), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[111]));   // sha_top.v(410)
    VERIFIC_DFFRS i3574 (.d(n2940), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[110]));   // sha_top.v(410)
    VERIFIC_DFFRS i3575 (.d(n2941), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[109]));   // sha_top.v(410)
    VERIFIC_DFFRS i3576 (.d(n2942), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[108]));   // sha_top.v(410)
    VERIFIC_DFFRS i3577 (.d(n2943), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[107]));   // sha_top.v(410)
    VERIFIC_DFFRS i3578 (.d(n2944), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[106]));   // sha_top.v(410)
    VERIFIC_DFFRS i3579 (.d(n2945), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[105]));   // sha_top.v(410)
    VERIFIC_DFFRS i3580 (.d(n2946), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[104]));   // sha_top.v(410)
    VERIFIC_DFFRS i3581 (.d(n2947), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[103]));   // sha_top.v(410)
    VERIFIC_DFFRS i3582 (.d(n2948), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[102]));   // sha_top.v(410)
    VERIFIC_DFFRS i3583 (.d(n2949), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[101]));   // sha_top.v(410)
    VERIFIC_DFFRS i3584 (.d(n2950), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[100]));   // sha_top.v(410)
    VERIFIC_DFFRS i3585 (.d(n2951), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[99]));   // sha_top.v(410)
    VERIFIC_DFFRS i3586 (.d(n2952), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[98]));   // sha_top.v(410)
    VERIFIC_DFFRS i3587 (.d(n2953), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[97]));   // sha_top.v(410)
    VERIFIC_DFFRS i3588 (.d(n2954), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[96]));   // sha_top.v(410)
    VERIFIC_DFFRS i3589 (.d(n2955), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[95]));   // sha_top.v(410)
    VERIFIC_DFFRS i3590 (.d(n2956), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[94]));   // sha_top.v(410)
    VERIFIC_DFFRS i3591 (.d(n2957), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[93]));   // sha_top.v(410)
    VERIFIC_DFFRS i3592 (.d(n2958), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[92]));   // sha_top.v(410)
    VERIFIC_DFFRS i3593 (.d(n2959), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[91]));   // sha_top.v(410)
    VERIFIC_DFFRS i3594 (.d(n2960), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[90]));   // sha_top.v(410)
    VERIFIC_DFFRS i3595 (.d(n2961), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[89]));   // sha_top.v(410)
    VERIFIC_DFFRS i3596 (.d(n2962), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[88]));   // sha_top.v(410)
    VERIFIC_DFFRS i3597 (.d(n2963), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[87]));   // sha_top.v(410)
    VERIFIC_DFFRS i3598 (.d(n2964), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[86]));   // sha_top.v(410)
    VERIFIC_DFFRS i3599 (.d(n2965), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[85]));   // sha_top.v(410)
    VERIFIC_DFFRS i3600 (.d(n2966), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[84]));   // sha_top.v(410)
    VERIFIC_DFFRS i3601 (.d(n2967), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[83]));   // sha_top.v(410)
    VERIFIC_DFFRS i3602 (.d(n2968), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[82]));   // sha_top.v(410)
    VERIFIC_DFFRS i3603 (.d(n2969), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[81]));   // sha_top.v(410)
    VERIFIC_DFFRS i3604 (.d(n2970), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[80]));   // sha_top.v(410)
    VERIFIC_DFFRS i3605 (.d(n2971), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[79]));   // sha_top.v(410)
    VERIFIC_DFFRS i3606 (.d(n2972), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[78]));   // sha_top.v(410)
    VERIFIC_DFFRS i3607 (.d(n2973), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[77]));   // sha_top.v(410)
    VERIFIC_DFFRS i3608 (.d(n2974), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[76]));   // sha_top.v(410)
    VERIFIC_DFFRS i3609 (.d(n2975), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[75]));   // sha_top.v(410)
    VERIFIC_DFFRS i3610 (.d(n2976), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[74]));   // sha_top.v(410)
    VERIFIC_DFFRS i3611 (.d(n2977), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[73]));   // sha_top.v(410)
    VERIFIC_DFFRS i3612 (.d(n2978), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[72]));   // sha_top.v(410)
    VERIFIC_DFFRS i3613 (.d(n2979), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[71]));   // sha_top.v(410)
    VERIFIC_DFFRS i3614 (.d(n2980), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[70]));   // sha_top.v(410)
    VERIFIC_DFFRS i3615 (.d(n2981), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[69]));   // sha_top.v(410)
    VERIFIC_DFFRS i3616 (.d(n2982), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[68]));   // sha_top.v(410)
    VERIFIC_DFFRS i3617 (.d(n2983), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[67]));   // sha_top.v(410)
    VERIFIC_DFFRS i3618 (.d(n2984), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[66]));   // sha_top.v(410)
    VERIFIC_DFFRS i3619 (.d(n2985), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[65]));   // sha_top.v(410)
    VERIFIC_DFFRS i3620 (.d(n2986), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[64]));   // sha_top.v(410)
    VERIFIC_DFFRS i3621 (.d(n2987), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[63]));   // sha_top.v(410)
    VERIFIC_DFFRS i3622 (.d(n2988), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[62]));   // sha_top.v(410)
    VERIFIC_DFFRS i3623 (.d(n2989), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[61]));   // sha_top.v(410)
    VERIFIC_DFFRS i3624 (.d(n2990), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[60]));   // sha_top.v(410)
    VERIFIC_DFFRS i3625 (.d(n2991), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[59]));   // sha_top.v(410)
    VERIFIC_DFFRS i3626 (.d(n2992), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[58]));   // sha_top.v(410)
    VERIFIC_DFFRS i3627 (.d(n2993), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[57]));   // sha_top.v(410)
    VERIFIC_DFFRS i3628 (.d(n2994), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[56]));   // sha_top.v(410)
    VERIFIC_DFFRS i3629 (.d(n2995), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[55]));   // sha_top.v(410)
    VERIFIC_DFFRS i3630 (.d(n2996), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[54]));   // sha_top.v(410)
    VERIFIC_DFFRS i3631 (.d(n2997), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[53]));   // sha_top.v(410)
    VERIFIC_DFFRS i3632 (.d(n2998), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[52]));   // sha_top.v(410)
    VERIFIC_DFFRS i3633 (.d(n2999), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[51]));   // sha_top.v(410)
    VERIFIC_DFFRS i3634 (.d(n3000), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[50]));   // sha_top.v(410)
    VERIFIC_DFFRS i3635 (.d(n3001), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[49]));   // sha_top.v(410)
    VERIFIC_DFFRS i3636 (.d(n3002), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[48]));   // sha_top.v(410)
    VERIFIC_DFFRS i3637 (.d(n3003), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[47]));   // sha_top.v(410)
    VERIFIC_DFFRS i3638 (.d(n3004), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[46]));   // sha_top.v(410)
    VERIFIC_DFFRS i3639 (.d(n3005), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[45]));   // sha_top.v(410)
    VERIFIC_DFFRS i3640 (.d(n3006), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[44]));   // sha_top.v(410)
    VERIFIC_DFFRS i3641 (.d(n3007), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[43]));   // sha_top.v(410)
    VERIFIC_DFFRS i3642 (.d(n3008), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[42]));   // sha_top.v(410)
    VERIFIC_DFFRS i3643 (.d(n3009), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[41]));   // sha_top.v(410)
    VERIFIC_DFFRS i3644 (.d(n3010), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[40]));   // sha_top.v(410)
    VERIFIC_DFFRS i3645 (.d(n3011), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[39]));   // sha_top.v(410)
    VERIFIC_DFFRS i3646 (.d(n3012), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[38]));   // sha_top.v(410)
    VERIFIC_DFFRS i3647 (.d(n3013), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[37]));   // sha_top.v(410)
    VERIFIC_DFFRS i3648 (.d(n3014), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[36]));   // sha_top.v(410)
    VERIFIC_DFFRS i3649 (.d(n3015), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[35]));   // sha_top.v(410)
    VERIFIC_DFFRS i3650 (.d(n3016), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[34]));   // sha_top.v(410)
    VERIFIC_DFFRS i3651 (.d(n3017), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[33]));   // sha_top.v(410)
    VERIFIC_DFFRS i3652 (.d(n3018), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[32]));   // sha_top.v(410)
    VERIFIC_DFFRS i3653 (.d(n3019), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[31]));   // sha_top.v(410)
    VERIFIC_DFFRS i3654 (.d(n3020), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[30]));   // sha_top.v(410)
    VERIFIC_DFFRS i3655 (.d(n3021), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[29]));   // sha_top.v(410)
    VERIFIC_DFFRS i3656 (.d(n3022), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[28]));   // sha_top.v(410)
    VERIFIC_DFFRS i3657 (.d(n3023), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[27]));   // sha_top.v(410)
    VERIFIC_DFFRS i3658 (.d(n3024), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[26]));   // sha_top.v(410)
    VERIFIC_DFFRS i3659 (.d(n3025), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[25]));   // sha_top.v(410)
    VERIFIC_DFFRS i3660 (.d(n3026), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[24]));   // sha_top.v(410)
    VERIFIC_DFFRS i3661 (.d(n3027), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[23]));   // sha_top.v(410)
    VERIFIC_DFFRS i3662 (.d(n3028), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[22]));   // sha_top.v(410)
    VERIFIC_DFFRS i3663 (.d(n3029), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[21]));   // sha_top.v(410)
    VERIFIC_DFFRS i3664 (.d(n3030), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[20]));   // sha_top.v(410)
    VERIFIC_DFFRS i3665 (.d(n3031), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[19]));   // sha_top.v(410)
    VERIFIC_DFFRS i3666 (.d(n3032), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[18]));   // sha_top.v(410)
    VERIFIC_DFFRS i3667 (.d(n3033), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[17]));   // sha_top.v(410)
    VERIFIC_DFFRS i3668 (.d(n3034), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[16]));   // sha_top.v(410)
    VERIFIC_DFFRS i3669 (.d(n3035), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[15]));   // sha_top.v(410)
    VERIFIC_DFFRS i3670 (.d(n3036), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[14]));   // sha_top.v(410)
    VERIFIC_DFFRS i3671 (.d(n3037), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[13]));   // sha_top.v(410)
    VERIFIC_DFFRS i3672 (.d(n3038), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[12]));   // sha_top.v(410)
    VERIFIC_DFFRS i3673 (.d(n3039), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[11]));   // sha_top.v(410)
    VERIFIC_DFFRS i3674 (.d(n3040), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[10]));   // sha_top.v(410)
    VERIFIC_DFFRS i3675 (.d(n3041), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[9]));   // sha_top.v(410)
    VERIFIC_DFFRS i3676 (.d(n3042), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[8]));   // sha_top.v(410)
    VERIFIC_DFFRS i3677 (.d(n3043), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[7]));   // sha_top.v(410)
    VERIFIC_DFFRS i3678 (.d(n3044), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[6]));   // sha_top.v(410)
    VERIFIC_DFFRS i3679 (.d(n3045), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[5]));   // sha_top.v(410)
    VERIFIC_DFFRS i3680 (.d(n3046), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[4]));   // sha_top.v(410)
    VERIFIC_DFFRS i3681 (.d(n3047), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[3]));   // sha_top.v(410)
    VERIFIC_DFFRS i3682 (.d(n3048), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[2]));   // sha_top.v(410)
    VERIFIC_DFFRS i3683 (.d(n3049), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3684 (.d(n3050), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_block[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3685 (.d(n3051), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[15]));   // sha_top.v(410)
    VERIFIC_DFFRS i3686 (.d(n3052), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[14]));   // sha_top.v(410)
    VERIFIC_DFFRS i3687 (.d(n3053), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[13]));   // sha_top.v(410)
    VERIFIC_DFFRS i3688 (.d(n3054), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[12]));   // sha_top.v(410)
    VERIFIC_DFFRS i3689 (.d(n3055), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[11]));   // sha_top.v(410)
    VERIFIC_DFFRS i3690 (.d(n3056), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[10]));   // sha_top.v(410)
    VERIFIC_DFFRS i3691 (.d(n3057), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[9]));   // sha_top.v(410)
    VERIFIC_DFFRS i3692 (.d(n3058), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[8]));   // sha_top.v(410)
    VERIFIC_DFFRS i3693 (.d(n3059), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[7]));   // sha_top.v(410)
    VERIFIC_DFFRS i3694 (.d(n3060), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[6]));   // sha_top.v(410)
    VERIFIC_DFFRS i3695 (.d(n3061), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[5]));   // sha_top.v(410)
    VERIFIC_DFFRS i3696 (.d(n3062), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[4]));   // sha_top.v(410)
    VERIFIC_DFFRS i3697 (.d(n3063), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[3]));   // sha_top.v(410)
    VERIFIC_DFFRS i3698 (.d(n3064), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[2]));   // sha_top.v(410)
    VERIFIC_DFFRS i3699 (.d(n3065), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3700 (.d(n3066), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_bytes_read[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3701 (.d(n3067), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[15]));   // sha_top.v(410)
    VERIFIC_DFFRS i3702 (.d(n3068), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[14]));   // sha_top.v(410)
    VERIFIC_DFFRS i3703 (.d(n3069), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[13]));   // sha_top.v(410)
    VERIFIC_DFFRS i3704 (.d(n3070), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[12]));   // sha_top.v(410)
    VERIFIC_DFFRS i3705 (.d(n3071), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[11]));   // sha_top.v(410)
    VERIFIC_DFFRS i3706 (.d(n3072), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[10]));   // sha_top.v(410)
    VERIFIC_DFFRS i3707 (.d(n3073), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[9]));   // sha_top.v(410)
    VERIFIC_DFFRS i3708 (.d(n3074), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[8]));   // sha_top.v(410)
    VERIFIC_DFFRS i3709 (.d(n3075), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[7]));   // sha_top.v(410)
    VERIFIC_DFFRS i3710 (.d(n3076), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[6]));   // sha_top.v(410)
    VERIFIC_DFFRS i3711 (.d(n3077), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[5]));   // sha_top.v(410)
    VERIFIC_DFFRS i3712 (.d(n3078), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[4]));   // sha_top.v(410)
    VERIFIC_DFFRS i3713 (.d(n3079), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[3]));   // sha_top.v(410)
    VERIFIC_DFFRS i3714 (.d(n3080), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[2]));   // sha_top.v(410)
    VERIFIC_DFFRS i3715 (.d(n3081), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3716 (.d(n3082), .clk(clk), .s(1'b0), .r(1'b0), .q(block_counter[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3717 (.d(n3083), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[159]));   // sha_top.v(410)
    VERIFIC_DFFRS i3718 (.d(n3084), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[158]));   // sha_top.v(410)
    VERIFIC_DFFRS i3719 (.d(n3085), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[157]));   // sha_top.v(410)
    VERIFIC_DFFRS i3720 (.d(n3086), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[156]));   // sha_top.v(410)
    VERIFIC_DFFRS i3721 (.d(n3087), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[155]));   // sha_top.v(410)
    VERIFIC_DFFRS i3722 (.d(n3088), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[154]));   // sha_top.v(410)
    VERIFIC_DFFRS i3723 (.d(n3089), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[153]));   // sha_top.v(410)
    VERIFIC_DFFRS i3724 (.d(n3090), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[152]));   // sha_top.v(410)
    VERIFIC_DFFRS i3725 (.d(n3091), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[151]));   // sha_top.v(410)
    VERIFIC_DFFRS i3726 (.d(n3092), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[150]));   // sha_top.v(410)
    VERIFIC_DFFRS i3727 (.d(n3093), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[149]));   // sha_top.v(410)
    VERIFIC_DFFRS i3728 (.d(n3094), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[148]));   // sha_top.v(410)
    VERIFIC_DFFRS i3729 (.d(n3095), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[147]));   // sha_top.v(410)
    VERIFIC_DFFRS i3730 (.d(n3096), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[146]));   // sha_top.v(410)
    VERIFIC_DFFRS i3731 (.d(n3097), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[145]));   // sha_top.v(410)
    VERIFIC_DFFRS i3732 (.d(n3098), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[144]));   // sha_top.v(410)
    VERIFIC_DFFRS i3733 (.d(n3099), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[143]));   // sha_top.v(410)
    VERIFIC_DFFRS i3734 (.d(n3100), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[142]));   // sha_top.v(410)
    VERIFIC_DFFRS i3735 (.d(n3101), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[141]));   // sha_top.v(410)
    VERIFIC_DFFRS i3736 (.d(n3102), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[140]));   // sha_top.v(410)
    VERIFIC_DFFRS i3737 (.d(n3103), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[139]));   // sha_top.v(410)
    VERIFIC_DFFRS i3738 (.d(n3104), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[138]));   // sha_top.v(410)
    VERIFIC_DFFRS i3739 (.d(n3105), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[137]));   // sha_top.v(410)
    VERIFIC_DFFRS i3740 (.d(n3106), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[136]));   // sha_top.v(410)
    VERIFIC_DFFRS i3741 (.d(n3107), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[135]));   // sha_top.v(410)
    VERIFIC_DFFRS i3742 (.d(n3108), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[134]));   // sha_top.v(410)
    VERIFIC_DFFRS i3743 (.d(n3109), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[133]));   // sha_top.v(410)
    VERIFIC_DFFRS i3744 (.d(n3110), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[132]));   // sha_top.v(410)
    VERIFIC_DFFRS i3745 (.d(n3111), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[131]));   // sha_top.v(410)
    VERIFIC_DFFRS i3746 (.d(n3112), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[130]));   // sha_top.v(410)
    VERIFIC_DFFRS i3747 (.d(n3113), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[129]));   // sha_top.v(410)
    VERIFIC_DFFRS i3748 (.d(n3114), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[128]));   // sha_top.v(410)
    VERIFIC_DFFRS i3749 (.d(n3115), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[127]));   // sha_top.v(410)
    VERIFIC_DFFRS i3750 (.d(n3116), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[126]));   // sha_top.v(410)
    VERIFIC_DFFRS i3751 (.d(n3117), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[125]));   // sha_top.v(410)
    VERIFIC_DFFRS i3752 (.d(n3118), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[124]));   // sha_top.v(410)
    VERIFIC_DFFRS i3753 (.d(n3119), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[123]));   // sha_top.v(410)
    VERIFIC_DFFRS i3754 (.d(n3120), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[122]));   // sha_top.v(410)
    VERIFIC_DFFRS i3755 (.d(n3121), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[121]));   // sha_top.v(410)
    VERIFIC_DFFRS i3756 (.d(n3122), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[120]));   // sha_top.v(410)
    VERIFIC_DFFRS i3757 (.d(n3123), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[119]));   // sha_top.v(410)
    VERIFIC_DFFRS i3758 (.d(n3124), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[118]));   // sha_top.v(410)
    VERIFIC_DFFRS i3759 (.d(n3125), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[117]));   // sha_top.v(410)
    VERIFIC_DFFRS i3760 (.d(n3126), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[116]));   // sha_top.v(410)
    VERIFIC_DFFRS i3761 (.d(n3127), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[115]));   // sha_top.v(410)
    VERIFIC_DFFRS i3762 (.d(n3128), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[114]));   // sha_top.v(410)
    VERIFIC_DFFRS i3763 (.d(n3129), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[113]));   // sha_top.v(410)
    VERIFIC_DFFRS i3764 (.d(n3130), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[112]));   // sha_top.v(410)
    VERIFIC_DFFRS i3765 (.d(n3131), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[111]));   // sha_top.v(410)
    VERIFIC_DFFRS i3766 (.d(n3132), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[110]));   // sha_top.v(410)
    VERIFIC_DFFRS i3767 (.d(n3133), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[109]));   // sha_top.v(410)
    VERIFIC_DFFRS i3768 (.d(n3134), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[108]));   // sha_top.v(410)
    VERIFIC_DFFRS i3769 (.d(n3135), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[107]));   // sha_top.v(410)
    VERIFIC_DFFRS i3770 (.d(n3136), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[106]));   // sha_top.v(410)
    VERIFIC_DFFRS i3771 (.d(n3137), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[105]));   // sha_top.v(410)
    VERIFIC_DFFRS i3772 (.d(n3138), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[104]));   // sha_top.v(410)
    VERIFIC_DFFRS i3773 (.d(n3139), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[103]));   // sha_top.v(410)
    VERIFIC_DFFRS i3774 (.d(n3140), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[102]));   // sha_top.v(410)
    VERIFIC_DFFRS i3775 (.d(n3141), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[101]));   // sha_top.v(410)
    VERIFIC_DFFRS i3776 (.d(n3142), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[100]));   // sha_top.v(410)
    VERIFIC_DFFRS i3777 (.d(n3143), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[99]));   // sha_top.v(410)
    VERIFIC_DFFRS i3778 (.d(n3144), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[98]));   // sha_top.v(410)
    VERIFIC_DFFRS i3779 (.d(n3145), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[97]));   // sha_top.v(410)
    VERIFIC_DFFRS i3780 (.d(n3146), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[96]));   // sha_top.v(410)
    VERIFIC_DFFRS i3781 (.d(n3147), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[95]));   // sha_top.v(410)
    VERIFIC_DFFRS i3782 (.d(n3148), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[94]));   // sha_top.v(410)
    VERIFIC_DFFRS i3783 (.d(n3149), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[93]));   // sha_top.v(410)
    VERIFIC_DFFRS i3784 (.d(n3150), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[92]));   // sha_top.v(410)
    VERIFIC_DFFRS i3785 (.d(n3151), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[91]));   // sha_top.v(410)
    VERIFIC_DFFRS i3786 (.d(n3152), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[90]));   // sha_top.v(410)
    VERIFIC_DFFRS i3787 (.d(n3153), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[89]));   // sha_top.v(410)
    VERIFIC_DFFRS i3788 (.d(n3154), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[88]));   // sha_top.v(410)
    VERIFIC_DFFRS i3789 (.d(n3155), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[87]));   // sha_top.v(410)
    VERIFIC_DFFRS i3790 (.d(n3156), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[86]));   // sha_top.v(410)
    VERIFIC_DFFRS i3791 (.d(n3157), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[85]));   // sha_top.v(410)
    VERIFIC_DFFRS i3792 (.d(n3158), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[84]));   // sha_top.v(410)
    VERIFIC_DFFRS i3793 (.d(n3159), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[83]));   // sha_top.v(410)
    VERIFIC_DFFRS i3794 (.d(n3160), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[82]));   // sha_top.v(410)
    VERIFIC_DFFRS i3795 (.d(n3161), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[81]));   // sha_top.v(410)
    VERIFIC_DFFRS i3796 (.d(n3162), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[80]));   // sha_top.v(410)
    VERIFIC_DFFRS i3797 (.d(n3163), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[79]));   // sha_top.v(410)
    VERIFIC_DFFRS i3798 (.d(n3164), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[78]));   // sha_top.v(410)
    VERIFIC_DFFRS i3799 (.d(n3165), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[77]));   // sha_top.v(410)
    VERIFIC_DFFRS i3800 (.d(n3166), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[76]));   // sha_top.v(410)
    VERIFIC_DFFRS i3801 (.d(n3167), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[75]));   // sha_top.v(410)
    VERIFIC_DFFRS i3802 (.d(n3168), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[74]));   // sha_top.v(410)
    VERIFIC_DFFRS i3803 (.d(n3169), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[73]));   // sha_top.v(410)
    VERIFIC_DFFRS i3804 (.d(n3170), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[72]));   // sha_top.v(410)
    VERIFIC_DFFRS i3805 (.d(n3171), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[71]));   // sha_top.v(410)
    VERIFIC_DFFRS i3806 (.d(n3172), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[70]));   // sha_top.v(410)
    VERIFIC_DFFRS i3807 (.d(n3173), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[69]));   // sha_top.v(410)
    VERIFIC_DFFRS i3808 (.d(n3174), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[68]));   // sha_top.v(410)
    VERIFIC_DFFRS i3809 (.d(n3175), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[67]));   // sha_top.v(410)
    VERIFIC_DFFRS i3810 (.d(n3176), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[66]));   // sha_top.v(410)
    VERIFIC_DFFRS i3811 (.d(n3177), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[65]));   // sha_top.v(410)
    VERIFIC_DFFRS i3812 (.d(n3178), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[64]));   // sha_top.v(410)
    VERIFIC_DFFRS i3813 (.d(n3179), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[63]));   // sha_top.v(410)
    VERIFIC_DFFRS i3814 (.d(n3180), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[62]));   // sha_top.v(410)
    VERIFIC_DFFRS i3815 (.d(n3181), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[61]));   // sha_top.v(410)
    VERIFIC_DFFRS i3816 (.d(n3182), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[60]));   // sha_top.v(410)
    VERIFIC_DFFRS i3817 (.d(n3183), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[59]));   // sha_top.v(410)
    VERIFIC_DFFRS i3818 (.d(n3184), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[58]));   // sha_top.v(410)
    VERIFIC_DFFRS i3819 (.d(n3185), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[57]));   // sha_top.v(410)
    VERIFIC_DFFRS i3820 (.d(n3186), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[56]));   // sha_top.v(410)
    VERIFIC_DFFRS i3821 (.d(n3187), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[55]));   // sha_top.v(410)
    VERIFIC_DFFRS i3822 (.d(n3188), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[54]));   // sha_top.v(410)
    VERIFIC_DFFRS i3823 (.d(n3189), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[53]));   // sha_top.v(410)
    VERIFIC_DFFRS i3824 (.d(n3190), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[52]));   // sha_top.v(410)
    VERIFIC_DFFRS i3825 (.d(n3191), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[51]));   // sha_top.v(410)
    VERIFIC_DFFRS i3826 (.d(n3192), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[50]));   // sha_top.v(410)
    VERIFIC_DFFRS i3827 (.d(n3193), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[49]));   // sha_top.v(410)
    VERIFIC_DFFRS i3828 (.d(n3194), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[48]));   // sha_top.v(410)
    VERIFIC_DFFRS i3829 (.d(n3195), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[47]));   // sha_top.v(410)
    VERIFIC_DFFRS i3830 (.d(n3196), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[46]));   // sha_top.v(410)
    VERIFIC_DFFRS i3831 (.d(n3197), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[45]));   // sha_top.v(410)
    VERIFIC_DFFRS i3832 (.d(n3198), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[44]));   // sha_top.v(410)
    VERIFIC_DFFRS i3833 (.d(n3199), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[43]));   // sha_top.v(410)
    VERIFIC_DFFRS i3834 (.d(n3200), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[42]));   // sha_top.v(410)
    VERIFIC_DFFRS i3835 (.d(n3201), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[41]));   // sha_top.v(410)
    VERIFIC_DFFRS i3836 (.d(n3202), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[40]));   // sha_top.v(410)
    VERIFIC_DFFRS i3837 (.d(n3203), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[39]));   // sha_top.v(410)
    VERIFIC_DFFRS i3838 (.d(n3204), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[38]));   // sha_top.v(410)
    VERIFIC_DFFRS i3839 (.d(n3205), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[37]));   // sha_top.v(410)
    VERIFIC_DFFRS i3840 (.d(n3206), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[36]));   // sha_top.v(410)
    VERIFIC_DFFRS i3841 (.d(n3207), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[35]));   // sha_top.v(410)
    VERIFIC_DFFRS i3842 (.d(n3208), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[34]));   // sha_top.v(410)
    VERIFIC_DFFRS i3843 (.d(n3209), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[33]));   // sha_top.v(410)
    VERIFIC_DFFRS i3844 (.d(n3210), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[32]));   // sha_top.v(410)
    VERIFIC_DFFRS i3845 (.d(n3211), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[31]));   // sha_top.v(410)
    VERIFIC_DFFRS i3846 (.d(n3212), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[30]));   // sha_top.v(410)
    VERIFIC_DFFRS i3847 (.d(n3213), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[29]));   // sha_top.v(410)
    VERIFIC_DFFRS i3848 (.d(n3214), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[28]));   // sha_top.v(410)
    VERIFIC_DFFRS i3849 (.d(n3215), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[27]));   // sha_top.v(410)
    VERIFIC_DFFRS i3850 (.d(n3216), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[26]));   // sha_top.v(410)
    VERIFIC_DFFRS i3851 (.d(n3217), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[25]));   // sha_top.v(410)
    VERIFIC_DFFRS i3852 (.d(n3218), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[24]));   // sha_top.v(410)
    VERIFIC_DFFRS i3853 (.d(n3219), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[23]));   // sha_top.v(410)
    VERIFIC_DFFRS i3854 (.d(n3220), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[22]));   // sha_top.v(410)
    VERIFIC_DFFRS i3855 (.d(n3221), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[21]));   // sha_top.v(410)
    VERIFIC_DFFRS i3856 (.d(n3222), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[20]));   // sha_top.v(410)
    VERIFIC_DFFRS i3857 (.d(n3223), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[19]));   // sha_top.v(410)
    VERIFIC_DFFRS i3858 (.d(n3224), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[18]));   // sha_top.v(410)
    VERIFIC_DFFRS i3859 (.d(n3225), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[17]));   // sha_top.v(410)
    VERIFIC_DFFRS i3860 (.d(n3226), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[16]));   // sha_top.v(410)
    VERIFIC_DFFRS i3861 (.d(n3227), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[15]));   // sha_top.v(410)
    VERIFIC_DFFRS i3862 (.d(n3228), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[14]));   // sha_top.v(410)
    VERIFIC_DFFRS i3863 (.d(n3229), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[13]));   // sha_top.v(410)
    VERIFIC_DFFRS i3864 (.d(n3230), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[12]));   // sha_top.v(410)
    VERIFIC_DFFRS i3865 (.d(n3231), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[11]));   // sha_top.v(410)
    VERIFIC_DFFRS i3866 (.d(n3232), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[10]));   // sha_top.v(410)
    VERIFIC_DFFRS i3867 (.d(n3233), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[9]));   // sha_top.v(410)
    VERIFIC_DFFRS i3868 (.d(n3234), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[8]));   // sha_top.v(410)
    VERIFIC_DFFRS i3869 (.d(n3235), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[7]));   // sha_top.v(410)
    VERIFIC_DFFRS i3870 (.d(n3236), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[6]));   // sha_top.v(410)
    VERIFIC_DFFRS i3871 (.d(n3237), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[5]));   // sha_top.v(410)
    VERIFIC_DFFRS i3872 (.d(n3238), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[4]));   // sha_top.v(410)
    VERIFIC_DFFRS i3873 (.d(n3239), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[3]));   // sha_top.v(410)
    VERIFIC_DFFRS i3874 (.d(n3240), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[2]));   // sha_top.v(410)
    VERIFIC_DFFRS i3875 (.d(n3241), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[1]));   // sha_top.v(410)
    VERIFIC_DFFRS i3876 (.d(n3242), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_reg_digest[0]));   // sha_top.v(410)
    VERIFIC_DFFRS i3877 (.d(n3243), .clk(clk), .s(1'b0), .r(1'b0), .q(sha_core_ready_r));   // sha_top.v(410)
    
endmodule

//
// Verific Verilog Description of OPERATOR LessThan_16u_16u
//

module LessThan_16u_16u (cin, a, b, o);
    input cin;
    input [15:0]a;
    input [15:0]b;
    output o;
    
    
    wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
        n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
        n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;
    
    xor (n1, a[0], b[0]) ;
    assign n2 = n1 ? b[0] : cin;
    xor (n3, a[1], b[1]) ;
    assign n4 = n3 ? b[1] : n2;
    xor (n5, a[2], b[2]) ;
    assign n6 = n5 ? b[2] : n4;
    xor (n7, a[3], b[3]) ;
    assign n8 = n7 ? b[3] : n6;
    xor (n9, a[4], b[4]) ;
    assign n10 = n9 ? b[4] : n8;
    xor (n11, a[5], b[5]) ;
    assign n12 = n11 ? b[5] : n10;
    xor (n13, a[6], b[6]) ;
    assign n14 = n13 ? b[6] : n12;
    xor (n15, a[7], b[7]) ;
    assign n16 = n15 ? b[7] : n14;
    xor (n17, a[8], b[8]) ;
    assign n18 = n17 ? b[8] : n16;
    xor (n19, a[9], b[9]) ;
    assign n20 = n19 ? b[9] : n18;
    xor (n21, a[10], b[10]) ;
    assign n22 = n21 ? b[10] : n20;
    xor (n23, a[11], b[11]) ;
    assign n24 = n23 ? b[11] : n22;
    xor (n25, a[12], b[12]) ;
    assign n26 = n25 ? b[12] : n24;
    xor (n27, a[13], b[13]) ;
    assign n28 = n27 ? b[13] : n26;
    xor (n29, a[14], b[14]) ;
    assign n30 = n29 ? b[14] : n28;
    xor (n31, a[15], b[15]) ;
    assign o = n31 ? b[15] : n30;
    
endmodule

//
// Verific Verilog Description of OPERATOR add_6u_6u
//

module add_6u_6u (cin, a, b, o, cout);
    input cin;
    input [5:0]a;
    input [5:0]b;
    output [5:0]o;
    output cout;
    
    
    wire n2, n4, n6, n8, n10;
    
    VERIFIC_FADD i1 (.cin(cin), .a(a[0]), .b(b[0]), .o(o[0]), .cout(n2));
    VERIFIC_FADD i2 (.cin(n2), .a(a[1]), .b(b[1]), .o(o[1]), .cout(n4));
    VERIFIC_FADD i3 (.cin(n4), .a(a[2]), .b(b[2]), .o(o[2]), .cout(n6));
    VERIFIC_FADD i4 (.cin(n6), .a(a[3]), .b(b[3]), .o(o[3]), .cout(n8));
    VERIFIC_FADD i5 (.cin(n8), .a(a[4]), .b(b[4]), .o(o[4]), .cout(n10));
    VERIFIC_FADD i6 (.cin(n10), .a(a[5]), .b(b[5]), .o(o[5]), .cout(cout));
    
endmodule

//
// Verific Verilog Description of OPERATOR add_16u_16u
//

module add_16u_16u (cin, a, b, o, cout);
    input cin;
    input [15:0]a;
    input [15:0]b;
    output [15:0]o;
    output cout;
    
    
    wire n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, 
        n24, n26, n28, n30;
    
    VERIFIC_FADD i1 (.cin(cin), .a(a[0]), .b(b[0]), .o(o[0]), .cout(n2));
    VERIFIC_FADD i2 (.cin(n2), .a(a[1]), .b(b[1]), .o(o[1]), .cout(n4));
    VERIFIC_FADD i3 (.cin(n4), .a(a[2]), .b(b[2]), .o(o[2]), .cout(n6));
    VERIFIC_FADD i4 (.cin(n6), .a(a[3]), .b(b[3]), .o(o[3]), .cout(n8));
    VERIFIC_FADD i5 (.cin(n8), .a(a[4]), .b(b[4]), .o(o[4]), .cout(n10));
    VERIFIC_FADD i6 (.cin(n10), .a(a[5]), .b(b[5]), .o(o[5]), .cout(n12));
    VERIFIC_FADD i7 (.cin(n12), .a(a[6]), .b(b[6]), .o(o[6]), .cout(n14));
    VERIFIC_FADD i8 (.cin(n14), .a(a[7]), .b(b[7]), .o(o[7]), .cout(n16));
    VERIFIC_FADD i9 (.cin(n16), .a(a[8]), .b(b[8]), .o(o[8]), .cout(n18));
    VERIFIC_FADD i10 (.cin(n18), .a(a[9]), .b(b[9]), .o(o[9]), .cout(n20));
    VERIFIC_FADD i11 (.cin(n20), .a(a[10]), .b(b[10]), .o(o[10]), .cout(n22));
    VERIFIC_FADD i12 (.cin(n22), .a(a[11]), .b(b[11]), .o(o[11]), .cout(n24));
    VERIFIC_FADD i13 (.cin(n24), .a(a[12]), .b(b[12]), .o(o[12]), .cout(n26));
    VERIFIC_FADD i14 (.cin(n26), .a(a[13]), .b(b[13]), .o(o[13]), .cout(n28));
    VERIFIC_FADD i15 (.cin(n28), .a(a[14]), .b(b[14]), .o(o[14]), .cout(n30));
    VERIFIC_FADD i16 (.cin(n30), .a(a[15]), .b(b[15]), .o(o[15]), .cout(cout));
    
endmodule

//
// Verific Verilog Description of OPERATOR add_10u_10u
//

module add_10u_10u (cin, a, b, o, cout);
    input cin;
    input [9:0]a;
    input [9:0]b;
    output [9:0]o;
    output cout;
    
    
    wire n2, n4, n6, n8, n10, n12, n14, n16, n18;
    
    VERIFIC_FADD i1 (.cin(cin), .a(a[0]), .b(b[0]), .o(o[0]), .cout(n2));
    VERIFIC_FADD i2 (.cin(n2), .a(a[1]), .b(b[1]), .o(o[1]), .cout(n4));
    VERIFIC_FADD i3 (.cin(n4), .a(a[2]), .b(b[2]), .o(o[2]), .cout(n6));
    VERIFIC_FADD i4 (.cin(n6), .a(a[3]), .b(b[3]), .o(o[3]), .cout(n8));
    VERIFIC_FADD i5 (.cin(n8), .a(a[4]), .b(b[4]), .o(o[4]), .cout(n10));
    VERIFIC_FADD i6 (.cin(n10), .a(a[5]), .b(b[5]), .o(o[5]), .cout(n12));
    VERIFIC_FADD i7 (.cin(n12), .a(a[6]), .b(b[6]), .o(o[6]), .cout(n14));
    VERIFIC_FADD i8 (.cin(n14), .a(a[7]), .b(b[7]), .o(o[7]), .cout(n16));
    VERIFIC_FADD i9 (.cin(n16), .a(a[8]), .b(b[8]), .o(o[8]), .cout(n18));
    VERIFIC_FADD i10 (.cin(n18), .a(a[9]), .b(b[9]), .o(o[9]), .cout(cout));
    
endmodule

//
// Verific Verilog Description of module reg2byte
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module sha1_core
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module modexp_top
//

module modexp_top (clk, rst, wr, addr, data_in, data_out, ack, 
            stb, in_addr_range, xram_addr, xram_data_out, xram_data_in, 
            xram_ack, xram_stb, xram_wr, exp_state, exp_addr, exp_step, 
            exp_m, exp_exp, exp_n, exp_valid);   // modexp_top.v(12)
    input clk;   // modexp_top.v(38)
    input rst;   // modexp_top.v(38)
    input wr;   // modexp_top.v(38)
    input [15:0]addr;   // modexp_top.v(40)
    input [7:0]data_in;   // modexp_top.v(39)
    output [7:0]data_out;   // modexp_top.v(41)
    output ack;   // modexp_top.v(42)
    input stb;   // modexp_top.v(38)
    output in_addr_range;   // modexp_top.v(43)
    output [15:0]xram_addr;   // modexp_top.v(46)
    output [7:0]xram_data_out;   // modexp_top.v(47)
    input [7:0]xram_data_in;   // modexp_top.v(48)
    input xram_ack;   // modexp_top.v(49)
    output xram_stb;   // modexp_top.v(50)
    output xram_wr;   // modexp_top.v(51)
    output [1:0]exp_state;   // modexp_top.v(54)
    output [15:0]exp_addr;   // modexp_top.v(55)
    output exp_step;   // modexp_top.v(57)
    output [2047:0]exp_m;   // modexp_top.v(56)
    output [2047:0]exp_exp;   // modexp_top.v(56)
    output [2047:0]exp_n;   // modexp_top.v(56)
    output exp_valid;   // modexp_top.v(57)
    
    wire sel_reg_start;   // modexp_top.v(84)
    wire sel_reg_state;   // modexp_top.v(85)
    wire sel_reg_addr;   // modexp_top.v(86)
    wire sel_reg_m;   // modexp_top.v(87)
    wire sel_reg_exp;   // modexp_top.v(88)
    wire sel_reg_n;   // modexp_top.v(89)
    wire exp_state_idle;   // modexp_top.v(103)
    wire exp_state_operate;   // modexp_top.v(104)
    wire exp_state_wait;   // modexp_top.v(105)
    wire wren;   // modexp_top.v(109)
    wire [7:0]exp_addr_dataout;   // modexp_top.v(114)
    wire [7:0]bigend_addr;   // modexp_top.v(128)
    wire [7:0]exp_m_dataout;   // modexp_top.v(132)
    wire [7:0]exp_exp_dataout;   // modexp_top.v(146)
    wire [7:0]exp_n_dataout;   // modexp_top.v(160)
    wire [7:0]byte_counter;   // modexp_top.v(179)
    wire reset_byte_counter;   // modexp_top.v(180)
    wire [7:0]byte_counter_next;   // modexp_top.v(182)
    wire last_byte_acked;   // modexp_top.v(186)
    wire [2:0]exp_reg_state_next_write_data;   // modexp_top.v(197)
    wire [2:0]exp_reg_state_next;   // modexp_top.v(199)
    wire [2047:0]exp_out;   // modexp_top.v(209)
    wire [2047:0]encrypted_data_buf;   // modexp_top.v(221)
    wire [2047:0]encrypted_data_buf_next;   // modexp_top.v(222)
    
    wire n4, n5, n8, n9, n10, n11, n12, n13, n14, n34, n56, 
        n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
        n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n97, n99, n105, n107, n116, n117, n118, n120, 
        n121, n122, n123, n124, n125, n126, n127, n129, n130, 
        n131, n132, n133, n134, n135, n136, n146, n147, n148, 
        n149, n150, n151, n152, n153, n176, n179, n180, n182, 
        n183, n187, n188, n2246, n2254, n2262, n2269, n2277, 
        n2284, n2291, n2297, n2305, n2312, n2319, n2325, n2332, 
        n2338, n2344, n2349, n2357, n2364, n2371, n2377, n2384, 
        n2390, n2396, n2401, n2408, n2414, n2420, n2425, n2431, 
        n2436, n2441, n2445, n2453, n2460, n2467, n2473, n2480, 
        n2486, n2492, n2497, n2504, n2510, n2516, n2521, n2527, 
        n2532, n2537, n2541, n2548, n2554, n2560, n2565, n2571, 
        n2576, n2581, n2585, n2591, n2596, n2601, n2605, n2610, 
        n2614, n2618, n2621, n2629, n2636, n2643, n2649, n2656, 
        n2662, n2668, n2673, n2680, n2686, n2692, n2697, n2703, 
        n2708, n2713, n2717, n2724, n2730, n2736, n2741, n2747, 
        n2752, n2757, n2761, n2767, n2772, n2777, n2781, n2786, 
        n2790, n2794, n2797, n2804, n2810, n2816, n2821, n2827, 
        n2832, n2837, n2841, n2847, n2852, n2857, n2861, n2866, 
        n2870, n2874, n2877, n2883, n2888, n2893, n2897, n2902, 
        n2906, n2910, n2913, n2918, n2922, n2926, n2929, n2933, 
        n2936, n2939, n2941, n2949, n2956, n2963, n2969, n2976, 
        n2982, n2988, n2993, n3000, n3006, n3012, n3017, n3023, 
        n3028, n3033, n3037, n3044, n3050, n3056, n3061, n3067, 
        n3072, n3077, n3081, n3087, n3092, n3097, n3101, n3106, 
        n3110, n3114, n3117, n3124, n3130, n3136, n3141, n3147, 
        n3152, n3157, n3161, n3167, n3172, n3177, n3181, n3186, 
        n3190, n3194, n3197, n3203, n3208, n3213, n3217, n3222, 
        n3226, n3230, n3233, n3238, n3242, n3246, n3249, n3253, 
        n3256, n3259, n3261, n3268, n3274, n3280, n3285, n3291, 
        n3296, n3301, n3305, n3311, n3316, n3321, n3325, n3330, 
        n3334, n3338, n3341, n3347, n3352, n3357, n3361, n3366, 
        n3370, n3374, n3377, n3382, n3386, n3390, n3393, n3397, 
        n3400, n3403, n3405, n3411, n3416, n3421, n3425, n3430, 
        n3434, n3438, n3441, n3446, n3450, n3454, n3457, n3461, 
        n3464, n3467, n3469, n3474, n3478, n3482, n3485, n3489, 
        n3492, n3495, n3497, n3501, n3504, n3507, n3509, n3512, 
        n3514, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
        n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, 
        n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
        n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
        n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, 
        n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
        n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, 
        n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
        n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
        n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
        n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
        n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, 
        n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
        n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
        n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, 
        n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
        n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, 
        n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
        n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, 
        n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, 
        n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
        n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, 
        n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
        n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, 
        n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
        n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
        n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, 
        n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
        n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, 
        n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, 
        n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
        n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, 
        n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, 
        n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, 
        n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, 
        n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
        n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, 
        n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
        n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, 
        n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, 
        n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
        n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
        n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
        n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, 
        n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
        n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
        n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
        n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
        n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
        n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, 
        n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
        n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
        n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
        n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
        n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, 
        n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
        n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, 
        n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
        n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
        n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
        n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
        n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
        n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
        n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
        n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
        n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
        n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, 
        n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
        n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
        n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
        n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
        n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
        n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
        n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
        n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, 
        n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
        n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, 
        n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
        n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
        n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
        n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
        n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, 
        n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
        n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
        n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, 
        n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
        n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, 
        n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
        n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
        n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
        n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
        n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, 
        n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
        n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
        n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
        n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
        n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
        n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
        n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
        n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
        n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
        n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, 
        n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
        n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, 
        n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
        n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
        n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
        n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
        n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
        n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
        n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
        n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
        n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
        n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
        n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
        n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
        n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, 
        n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
        n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, 
        n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
        n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
        n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
        n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
        n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
        n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
        n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
        n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
        n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
        n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
        n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
        n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
        n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
        n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
        n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
        n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
        n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
        n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
        n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
        n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
        n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, 
        n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
        n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
        n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
        n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
        n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, 
        n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
        n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, 
        n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, 
        n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
        n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, 
        n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
        n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, 
        n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
        n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, 
        n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, 
        n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
        n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, 
        n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
        n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
        n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, 
        n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
        n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, 
        n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, 
        n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
        n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, 
        n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
        n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, 
        n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
        n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, 
        n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, 
        n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
        n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, 
        n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, 
        n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, 
        n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, 
        n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
        n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
        n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, 
        n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, 
        n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, 
        n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
        n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, 
        n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, 
        n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, 
        n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, 
        n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
        n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
        n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, 
        n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, 
        n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, 
        n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
        n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, 
        n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, 
        n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, 
        n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, 
        n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
        n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
        n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, 
        n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, 
        n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, 
        n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
        n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, 
        n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, 
        n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, 
        n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, 
        n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
        n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, 
        n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, 
        n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, 
        n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, 
        n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
        n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, 
        n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, 
        n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, 
        n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, 
        n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, 
        n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, 
        n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, 
        n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, 
        n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
        n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
        n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, 
        n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, 
        n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, 
        n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
        n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
        n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, 
        n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, 
        n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, 
        n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
        n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
        n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, 
        n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, 
        n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, 
        n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, 
        n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
        n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, 
        n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, 
        n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, 
        n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, 
        n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, 
        n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, 
        n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, 
        n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, 
        n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, 
        n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
        n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, 
        n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, 
        n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, 
        n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
        n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
        n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, 
        n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, 
        n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, 
        n5547, n5548, n7616, n7617, n7618, n7619, n7620, n7621, 
        n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, 
        n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, 
        n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, 
        n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
        n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
        n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, 
        n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, 
        n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, 
        n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
        n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, 
        n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, 
        n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, 
        n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, 
        n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
        n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, 
        n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, 
        n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, 
        n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, 
        n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
        n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, 
        n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, 
        n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, 
        n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, 
        n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
        n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
        n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, 
        n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, 
        n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, 
        n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
        n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, 
        n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, 
        n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, 
        n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
        n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
        n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, 
        n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, 
        n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, 
        n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, 
        n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
        n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, 
        n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, 
        n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, 
        n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, 
        n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
        n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, 
        n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, 
        n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, 
        n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
        n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
        n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, 
        n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, 
        n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, 
        n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
        n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
        n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, 
        n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, 
        n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, 
        n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
        n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
        n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, 
        n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, 
        n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, 
        n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, 
        n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
        n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, 
        n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, 
        n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, 
        n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, 
        n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
        n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, 
        n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, 
        n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, 
        n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, 
        n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
        n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, 
        n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, 
        n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, 
        n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, 
        n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
        n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, 
        n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, 
        n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, 
        n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, 
        n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
        n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, 
        n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, 
        n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, 
        n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, 
        n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
        n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, 
        n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, 
        n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, 
        n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, 
        n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
        n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, 
        n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, 
        n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, 
        n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, 
        n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
        n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, 
        n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, 
        n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, 
        n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, 
        n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
        n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, 
        n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, 
        n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, 
        n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
        n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
        n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, 
        n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, 
        n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
        n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, 
        n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
        n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, 
        n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, 
        n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, 
        n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
        n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
        n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, 
        n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, 
        n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
        n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, 
        n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
        n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, 
        n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, 
        n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, 
        n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, 
        n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
        n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, 
        n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, 
        n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, 
        n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, 
        n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
        n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, 
        n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, 
        n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
        n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, 
        n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
        n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, 
        n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, 
        n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, 
        n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
        n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
        n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, 
        n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, 
        n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, 
        n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
        n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
        n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, 
        n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, 
        n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, 
        n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
        n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
        n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, 
        n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, 
        n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
        n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
        n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
        n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, 
        n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, 
        n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, 
        n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
        n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
        n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, 
        n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, 
        n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, 
        n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
        n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
        n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, 
        n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, 
        n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, 
        n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
        n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
        n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, 
        n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, 
        n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, 
        n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
        n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
        n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, 
        n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, 
        n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, 
        n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
        n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
        n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, 
        n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, 
        n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
        n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
        n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
        n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, 
        n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, 
        n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
        n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, 
        n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
        n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, 
        n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, 
        n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
        n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, 
        n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
        n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, 
        n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, 
        n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, 
        n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, 
        n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
        n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, 
        n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, 
        n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, 
        n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, 
        n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
        n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, 
        n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, 
        n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, 
        n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
        n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
        n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, 
        n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, 
        n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, 
        n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
        n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
        n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, 
        n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, 
        n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, 
        n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, 
        n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
        n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, 
        n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, 
        n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, 
        n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, 
        n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
        n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, 
        n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, 
        n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
        n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, 
        n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
        n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, 
        n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, 
        n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, 
        n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
        n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
        n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, 
        n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, 
        n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, 
        n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
        n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
        n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, 
        n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, 
        n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, 
        n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, 
        n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
        n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, 
        n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, 
        n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, 
        n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, 
        n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
        n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, 
        n9662, n9663;
    
    assign xram_stb = xram_wr;   // modexp_top.v(50)
    LessThan_16u_16u LessThan_3 (.cin(1'b1), .a({16'b1111101000000000}), 
            .b({addr}), .o(n4));   // modexp_top.v(81)
    LessThan_16u_16u LessThan_4 (.cin(1'b0), .a({addr}), .b({16'b1111110100010000}), 
            .o(n5));   // modexp_top.v(81)
    and (in_addr_range, n4, n5) ;   // modexp_top.v(81)
    and (ack, stb, in_addr_range) ;   // modexp_top.v(82)
    not (n8, addr[8]) ;   // modexp_top.v(84)
    not (n9, addr[10]) ;   // modexp_top.v(84)
    not (n10, addr[11]) ;   // modexp_top.v(84)
    not (n11, addr[12]) ;   // modexp_top.v(84)
    not (n12, addr[13]) ;   // modexp_top.v(84)
    not (n13, addr[14]) ;   // modexp_top.v(84)
    not (n14, addr[15]) ;   // modexp_top.v(84)
    nor (sel_reg_start, n14, n13, n12, n11, n10, n9, addr[9], 
        n8, addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], 
        addr[1], addr[0]) ;   // modexp_top.v(84)
    not (bigend_addr[0], addr[0]) ;   // modexp_top.v(85)
    nor (sel_reg_state, n14, n13, n12, n11, n10, n9, addr[9], 
        n8, addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], 
        addr[1], bigend_addr[0]) ;   // modexp_top.v(85)
    not (bigend_addr[1], addr[1]) ;   // modexp_top.v(86)
    nor (sel_reg_addr, n14, n13, n12, n11, n10, n9, addr[9], 
        n8, addr[7], addr[6], addr[5], addr[4], addr[3], addr[2], 
        bigend_addr[1]) ;   // modexp_top.v(86)
    not (n34, addr[9]) ;   // modexp_top.v(87)
    nor (sel_reg_m, n14, n13, n12, n11, n10, addr[10], n34, 
        addr[8]) ;   // modexp_top.v(87)
    nor (sel_reg_exp, n14, n13, n12, n11, n10, addr[10], n34, 
        n8) ;   // modexp_top.v(88)
    nor (sel_reg_n, n14, n13, n12, n11, n10, n9, addr[9], addr[8]) ;   // modexp_top.v(89)
    assign n56 = sel_reg_n ? exp_n_dataout[7] : 1'b0;   // modexp_top.v(100)
    assign n57 = sel_reg_n ? exp_n_dataout[6] : 1'b0;   // modexp_top.v(100)
    assign n58 = sel_reg_n ? exp_n_dataout[5] : 1'b0;   // modexp_top.v(100)
    assign n59 = sel_reg_n ? exp_n_dataout[4] : 1'b0;   // modexp_top.v(100)
    assign n60 = sel_reg_n ? exp_n_dataout[3] : 1'b0;   // modexp_top.v(100)
    assign n61 = sel_reg_n ? exp_n_dataout[2] : 1'b0;   // modexp_top.v(100)
    assign n62 = sel_reg_n ? exp_n_dataout[1] : 1'b0;   // modexp_top.v(100)
    assign n63 = sel_reg_n ? exp_n_dataout[0] : 1'b0;   // modexp_top.v(100)
    assign n64 = sel_reg_exp ? exp_exp_dataout[7] : n56;   // modexp_top.v(100)
    assign n65 = sel_reg_exp ? exp_exp_dataout[6] : n57;   // modexp_top.v(100)
    assign n66 = sel_reg_exp ? exp_exp_dataout[5] : n58;   // modexp_top.v(100)
    assign n67 = sel_reg_exp ? exp_exp_dataout[4] : n59;   // modexp_top.v(100)
    assign n68 = sel_reg_exp ? exp_exp_dataout[3] : n60;   // modexp_top.v(100)
    assign n69 = sel_reg_exp ? exp_exp_dataout[2] : n61;   // modexp_top.v(100)
    assign n70 = sel_reg_exp ? exp_exp_dataout[1] : n62;   // modexp_top.v(100)
    assign n71 = sel_reg_exp ? exp_exp_dataout[0] : n63;   // modexp_top.v(100)
    assign n72 = sel_reg_m ? exp_m_dataout[7] : n64;   // modexp_top.v(100)
    assign n73 = sel_reg_m ? exp_m_dataout[6] : n65;   // modexp_top.v(100)
    assign n74 = sel_reg_m ? exp_m_dataout[5] : n66;   // modexp_top.v(100)
    assign n75 = sel_reg_m ? exp_m_dataout[4] : n67;   // modexp_top.v(100)
    assign n76 = sel_reg_m ? exp_m_dataout[3] : n68;   // modexp_top.v(100)
    assign n77 = sel_reg_m ? exp_m_dataout[2] : n69;   // modexp_top.v(100)
    assign n78 = sel_reg_m ? exp_m_dataout[1] : n70;   // modexp_top.v(100)
    assign n79 = sel_reg_m ? exp_m_dataout[0] : n71;   // modexp_top.v(100)
    assign n80 = sel_reg_addr ? exp_addr_dataout[7] : n72;   // modexp_top.v(100)
    assign n81 = sel_reg_addr ? exp_addr_dataout[6] : n73;   // modexp_top.v(100)
    assign n82 = sel_reg_addr ? exp_addr_dataout[5] : n74;   // modexp_top.v(100)
    assign n83 = sel_reg_addr ? exp_addr_dataout[4] : n75;   // modexp_top.v(100)
    assign n84 = sel_reg_addr ? exp_addr_dataout[3] : n76;   // modexp_top.v(100)
    assign n85 = sel_reg_addr ? exp_addr_dataout[2] : n77;   // modexp_top.v(100)
    assign n86 = sel_reg_addr ? exp_addr_dataout[1] : n78;   // modexp_top.v(100)
    assign n87 = sel_reg_addr ? exp_addr_dataout[0] : n79;   // modexp_top.v(100)
    assign data_out[7] = sel_reg_state ? 1'b0 : n80;   // modexp_top.v(100)
    assign data_out[6] = sel_reg_state ? 1'b0 : n81;   // modexp_top.v(100)
    assign data_out[5] = sel_reg_state ? 1'b0 : n82;   // modexp_top.v(100)
    assign data_out[4] = sel_reg_state ? 1'b0 : n83;   // modexp_top.v(100)
    assign data_out[3] = sel_reg_state ? 1'b0 : n84;   // modexp_top.v(100)
    assign data_out[2] = sel_reg_state ? 1'b0 : n85;   // modexp_top.v(100)
    assign data_out[1] = sel_reg_state ? exp_state[1] : n86;   // modexp_top.v(100)
    assign data_out[0] = sel_reg_state ? exp_state[0] : n87;   // modexp_top.v(100)
    nor (exp_state_idle, exp_state[1], exp_state[0]) ;   // modexp_top.v(103)
    not (n97, exp_state[0]) ;   // modexp_top.v(104)
    nor (exp_state_operate, exp_state[1], n97) ;   // modexp_top.v(104)
    not (n99, exp_state[1]) ;   // modexp_top.v(105)
    nor (exp_state_wait, n99, exp_state[0]) ;   // modexp_top.v(105)
    nor (xram_wr, n99, n97) ;   // modexp_top.v(106)
    and (wren, wr, exp_state_idle) ;   // modexp_top.v(109)
    and (n105, sel_reg_start, data_in[0]) ;   // modexp_top.v(110)
    and (reset_byte_counter, n105, wren) ;   // modexp_top.v(110)
    reg2byte exp_reg_opaddr_i (.clk(clk), .rst(rst), .en(sel_reg_addr), 
            .wr(n107), .addr(addr[0]), .data_in({data_in}), .data_out({exp_addr_dataout}), 
            .reg_out({exp_addr}));   // modexp_top.v(115)
    and (n107, sel_reg_addr, wren) ;   // modexp_top.v(119)
    not (bigend_addr[7], addr[7]) ;   // modexp_top.v(128)
    not (bigend_addr[6], addr[6]) ;   // modexp_top.v(128)
    not (bigend_addr[5], addr[5]) ;   // modexp_top.v(128)
    not (bigend_addr[4], addr[4]) ;   // modexp_top.v(128)
    not (bigend_addr[3], addr[3]) ;   // modexp_top.v(128)
    not (bigend_addr[2], addr[2]) ;   // modexp_top.v(128)
    reg256byte exp_reg_m_i (.clk(clk), .rst(rst), .en(sel_reg_m), .wr(n116), 
            .addr({bigend_addr}), .data_in({data_in}), .data_out({exp_m_dataout}), 
            .reg_out({exp_m}));   // modexp_top.v(133)
    and (n116, sel_reg_m, wren) ;   // modexp_top.v(137)
    reg256byte exp_reg_exp_i (.clk(clk), .rst(rst), .en(sel_reg_exp), 
            .wr(n117), .addr({bigend_addr}), .data_in({data_in}), .data_out({exp_exp_dataout}), 
            .reg_out({exp_exp}));   // modexp_top.v(147)
    and (n117, sel_reg_exp, wren) ;   // modexp_top.v(151)
    reg256byte exp_reg_n_i (.clk(clk), .rst(rst), .en(sel_reg_n), .wr(n118), 
            .addr({bigend_addr}), .data_in({data_in}), .data_out({exp_n_dataout}), 
            .reg_out({exp_n}));   // modexp_top.v(161)
    and (n118, sel_reg_n, wren) ;   // modexp_top.v(165)
    add_8u_8u add_118 (.cin(1'b0), .a({byte_counter}), .b({8'b00000001}), 
            .o({n120, n121, n122, n123, n124, n125, n126, n127}));   // modexp_top.v(183)
    assign n129 = xram_ack ? n120 : byte_counter[7];   // modexp_top.v(184)
    assign n130 = xram_ack ? n121 : byte_counter[6];   // modexp_top.v(184)
    assign n131 = xram_ack ? n122 : byte_counter[5];   // modexp_top.v(184)
    assign n132 = xram_ack ? n123 : byte_counter[4];   // modexp_top.v(184)
    assign n133 = xram_ack ? n124 : byte_counter[3];   // modexp_top.v(184)
    assign n134 = xram_ack ? n125 : byte_counter[2];   // modexp_top.v(184)
    assign n135 = xram_ack ? n126 : byte_counter[1];   // modexp_top.v(184)
    assign n136 = xram_ack ? n127 : byte_counter[0];   // modexp_top.v(184)
    assign byte_counter_next[7] = reset_byte_counter ? 1'b0 : n129;   // modexp_top.v(184)
    assign byte_counter_next[6] = reset_byte_counter ? 1'b0 : n130;   // modexp_top.v(184)
    assign byte_counter_next[5] = reset_byte_counter ? 1'b0 : n131;   // modexp_top.v(184)
    assign byte_counter_next[4] = reset_byte_counter ? 1'b0 : n132;   // modexp_top.v(184)
    assign byte_counter_next[3] = reset_byte_counter ? 1'b0 : n133;   // modexp_top.v(184)
    assign byte_counter_next[2] = reset_byte_counter ? 1'b0 : n134;   // modexp_top.v(184)
    assign byte_counter_next[1] = reset_byte_counter ? 1'b0 : n135;   // modexp_top.v(184)
    assign byte_counter_next[0] = reset_byte_counter ? 1'b0 : n136;   // modexp_top.v(184)
    not (n146, byte_counter[0]) ;   // modexp_top.v(186)
    not (n147, byte_counter[1]) ;   // modexp_top.v(186)
    not (n148, byte_counter[2]) ;   // modexp_top.v(186)
    not (n149, byte_counter[3]) ;   // modexp_top.v(186)
    not (n150, byte_counter[4]) ;   // modexp_top.v(186)
    not (n151, byte_counter[5]) ;   // modexp_top.v(186)
    not (n152, byte_counter[6]) ;   // modexp_top.v(186)
    not (n153, byte_counter[7]) ;   // modexp_top.v(186)
    nor (n2246, n153, n152, n151, n150, n149, n148, n147, n146) ;   // modexp_top.v(186)
    and (last_byte_acked, n2246, xram_ack) ;   // modexp_top.v(186)
    add_16u_16u add_147 (.cin(1'b0), .a({exp_addr}), .b({8'b00000000, 
            byte_counter}), .o({xram_addr}));   // modexp_top.v(189)
    not (exp_reg_state_next_write_data[1], last_byte_acked) ;   // modexp_top.v(197)
    assign n176 = xram_wr ? exp_reg_state_next_write_data[1] : 1'b0;   // modexp_top.v(204)
    assign n179 = exp_state_wait ? 1'b1 : n176;   // modexp_top.v(204)
    assign n180 = exp_state_wait ? exp_valid : n176;   // modexp_top.v(204)
    assign n182 = exp_state_operate ? 1'b1 : n179;   // modexp_top.v(204)
    assign n183 = exp_state_operate ? 1'b0 : n180;   // modexp_top.v(204)
    assign exp_reg_state_next[1] = exp_state_idle ? 1'b0 : n182;   // modexp_top.v(204)
    assign exp_reg_state_next[0] = exp_state_idle ? reset_byte_counter : n183;   // modexp_top.v(204)
    xor (n187, exp_state[0], exp_reg_state_next[0]) ;   // modexp_top.v(206)
    xor (n188, exp_state[1], exp_reg_state_next[1]) ;   // modexp_top.v(206)
    or (exp_step, n188, n187) ;   // modexp_top.v(206)
    modexp modexp_i (.clk(clk), .rst(rst), .start(reset_byte_counter), 
           .ready(exp_valid), .m({exp_m}), .e({exp_exp}), .n({exp_n}), 
           .c({exp_out}));   // modexp_top.v(210)
    assign encrypted_data_buf_next[2047] = exp_valid ? exp_out[2047] : encrypted_data_buf[2047];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2046] = exp_valid ? exp_out[2046] : encrypted_data_buf[2046];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2045] = exp_valid ? exp_out[2045] : encrypted_data_buf[2045];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2044] = exp_valid ? exp_out[2044] : encrypted_data_buf[2044];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2043] = exp_valid ? exp_out[2043] : encrypted_data_buf[2043];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2042] = exp_valid ? exp_out[2042] : encrypted_data_buf[2042];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2041] = exp_valid ? exp_out[2041] : encrypted_data_buf[2041];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2040] = exp_valid ? exp_out[2040] : encrypted_data_buf[2040];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2039] = exp_valid ? exp_out[2039] : encrypted_data_buf[2039];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2038] = exp_valid ? exp_out[2038] : encrypted_data_buf[2038];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2037] = exp_valid ? exp_out[2037] : encrypted_data_buf[2037];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2036] = exp_valid ? exp_out[2036] : encrypted_data_buf[2036];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2035] = exp_valid ? exp_out[2035] : encrypted_data_buf[2035];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2034] = exp_valid ? exp_out[2034] : encrypted_data_buf[2034];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2033] = exp_valid ? exp_out[2033] : encrypted_data_buf[2033];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2032] = exp_valid ? exp_out[2032] : encrypted_data_buf[2032];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2031] = exp_valid ? exp_out[2031] : encrypted_data_buf[2031];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2030] = exp_valid ? exp_out[2030] : encrypted_data_buf[2030];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2029] = exp_valid ? exp_out[2029] : encrypted_data_buf[2029];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2028] = exp_valid ? exp_out[2028] : encrypted_data_buf[2028];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2027] = exp_valid ? exp_out[2027] : encrypted_data_buf[2027];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2026] = exp_valid ? exp_out[2026] : encrypted_data_buf[2026];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2025] = exp_valid ? exp_out[2025] : encrypted_data_buf[2025];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2024] = exp_valid ? exp_out[2024] : encrypted_data_buf[2024];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2023] = exp_valid ? exp_out[2023] : encrypted_data_buf[2023];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2022] = exp_valid ? exp_out[2022] : encrypted_data_buf[2022];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2021] = exp_valid ? exp_out[2021] : encrypted_data_buf[2021];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2020] = exp_valid ? exp_out[2020] : encrypted_data_buf[2020];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2019] = exp_valid ? exp_out[2019] : encrypted_data_buf[2019];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2018] = exp_valid ? exp_out[2018] : encrypted_data_buf[2018];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2017] = exp_valid ? exp_out[2017] : encrypted_data_buf[2017];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2016] = exp_valid ? exp_out[2016] : encrypted_data_buf[2016];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2015] = exp_valid ? exp_out[2015] : encrypted_data_buf[2015];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2014] = exp_valid ? exp_out[2014] : encrypted_data_buf[2014];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2013] = exp_valid ? exp_out[2013] : encrypted_data_buf[2013];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2012] = exp_valid ? exp_out[2012] : encrypted_data_buf[2012];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2011] = exp_valid ? exp_out[2011] : encrypted_data_buf[2011];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2010] = exp_valid ? exp_out[2010] : encrypted_data_buf[2010];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2009] = exp_valid ? exp_out[2009] : encrypted_data_buf[2009];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2008] = exp_valid ? exp_out[2008] : encrypted_data_buf[2008];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2007] = exp_valid ? exp_out[2007] : encrypted_data_buf[2007];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2006] = exp_valid ? exp_out[2006] : encrypted_data_buf[2006];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2005] = exp_valid ? exp_out[2005] : encrypted_data_buf[2005];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2004] = exp_valid ? exp_out[2004] : encrypted_data_buf[2004];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2003] = exp_valid ? exp_out[2003] : encrypted_data_buf[2003];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2002] = exp_valid ? exp_out[2002] : encrypted_data_buf[2002];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2001] = exp_valid ? exp_out[2001] : encrypted_data_buf[2001];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2000] = exp_valid ? exp_out[2000] : encrypted_data_buf[2000];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1999] = exp_valid ? exp_out[1999] : encrypted_data_buf[1999];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1998] = exp_valid ? exp_out[1998] : encrypted_data_buf[1998];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1997] = exp_valid ? exp_out[1997] : encrypted_data_buf[1997];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1996] = exp_valid ? exp_out[1996] : encrypted_data_buf[1996];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1995] = exp_valid ? exp_out[1995] : encrypted_data_buf[1995];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1994] = exp_valid ? exp_out[1994] : encrypted_data_buf[1994];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1993] = exp_valid ? exp_out[1993] : encrypted_data_buf[1993];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1992] = exp_valid ? exp_out[1992] : encrypted_data_buf[1992];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1991] = exp_valid ? exp_out[1991] : encrypted_data_buf[1991];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1990] = exp_valid ? exp_out[1990] : encrypted_data_buf[1990];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1989] = exp_valid ? exp_out[1989] : encrypted_data_buf[1989];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1988] = exp_valid ? exp_out[1988] : encrypted_data_buf[1988];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1987] = exp_valid ? exp_out[1987] : encrypted_data_buf[1987];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1986] = exp_valid ? exp_out[1986] : encrypted_data_buf[1986];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1985] = exp_valid ? exp_out[1985] : encrypted_data_buf[1985];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1984] = exp_valid ? exp_out[1984] : encrypted_data_buf[1984];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1983] = exp_valid ? exp_out[1983] : encrypted_data_buf[1983];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1982] = exp_valid ? exp_out[1982] : encrypted_data_buf[1982];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1981] = exp_valid ? exp_out[1981] : encrypted_data_buf[1981];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1980] = exp_valid ? exp_out[1980] : encrypted_data_buf[1980];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1979] = exp_valid ? exp_out[1979] : encrypted_data_buf[1979];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1978] = exp_valid ? exp_out[1978] : encrypted_data_buf[1978];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1977] = exp_valid ? exp_out[1977] : encrypted_data_buf[1977];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1976] = exp_valid ? exp_out[1976] : encrypted_data_buf[1976];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1975] = exp_valid ? exp_out[1975] : encrypted_data_buf[1975];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1974] = exp_valid ? exp_out[1974] : encrypted_data_buf[1974];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1973] = exp_valid ? exp_out[1973] : encrypted_data_buf[1973];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1972] = exp_valid ? exp_out[1972] : encrypted_data_buf[1972];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1971] = exp_valid ? exp_out[1971] : encrypted_data_buf[1971];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1970] = exp_valid ? exp_out[1970] : encrypted_data_buf[1970];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1969] = exp_valid ? exp_out[1969] : encrypted_data_buf[1969];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1968] = exp_valid ? exp_out[1968] : encrypted_data_buf[1968];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1967] = exp_valid ? exp_out[1967] : encrypted_data_buf[1967];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1966] = exp_valid ? exp_out[1966] : encrypted_data_buf[1966];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1965] = exp_valid ? exp_out[1965] : encrypted_data_buf[1965];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1964] = exp_valid ? exp_out[1964] : encrypted_data_buf[1964];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1963] = exp_valid ? exp_out[1963] : encrypted_data_buf[1963];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1962] = exp_valid ? exp_out[1962] : encrypted_data_buf[1962];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1961] = exp_valid ? exp_out[1961] : encrypted_data_buf[1961];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1960] = exp_valid ? exp_out[1960] : encrypted_data_buf[1960];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1959] = exp_valid ? exp_out[1959] : encrypted_data_buf[1959];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1958] = exp_valid ? exp_out[1958] : encrypted_data_buf[1958];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1957] = exp_valid ? exp_out[1957] : encrypted_data_buf[1957];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1956] = exp_valid ? exp_out[1956] : encrypted_data_buf[1956];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1955] = exp_valid ? exp_out[1955] : encrypted_data_buf[1955];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1954] = exp_valid ? exp_out[1954] : encrypted_data_buf[1954];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1953] = exp_valid ? exp_out[1953] : encrypted_data_buf[1953];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1952] = exp_valid ? exp_out[1952] : encrypted_data_buf[1952];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1951] = exp_valid ? exp_out[1951] : encrypted_data_buf[1951];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1950] = exp_valid ? exp_out[1950] : encrypted_data_buf[1950];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1949] = exp_valid ? exp_out[1949] : encrypted_data_buf[1949];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1948] = exp_valid ? exp_out[1948] : encrypted_data_buf[1948];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1947] = exp_valid ? exp_out[1947] : encrypted_data_buf[1947];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1946] = exp_valid ? exp_out[1946] : encrypted_data_buf[1946];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1945] = exp_valid ? exp_out[1945] : encrypted_data_buf[1945];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1944] = exp_valid ? exp_out[1944] : encrypted_data_buf[1944];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1943] = exp_valid ? exp_out[1943] : encrypted_data_buf[1943];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1942] = exp_valid ? exp_out[1942] : encrypted_data_buf[1942];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1941] = exp_valid ? exp_out[1941] : encrypted_data_buf[1941];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1940] = exp_valid ? exp_out[1940] : encrypted_data_buf[1940];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1939] = exp_valid ? exp_out[1939] : encrypted_data_buf[1939];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1938] = exp_valid ? exp_out[1938] : encrypted_data_buf[1938];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1937] = exp_valid ? exp_out[1937] : encrypted_data_buf[1937];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1936] = exp_valid ? exp_out[1936] : encrypted_data_buf[1936];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1935] = exp_valid ? exp_out[1935] : encrypted_data_buf[1935];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1934] = exp_valid ? exp_out[1934] : encrypted_data_buf[1934];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1933] = exp_valid ? exp_out[1933] : encrypted_data_buf[1933];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1932] = exp_valid ? exp_out[1932] : encrypted_data_buf[1932];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1931] = exp_valid ? exp_out[1931] : encrypted_data_buf[1931];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1930] = exp_valid ? exp_out[1930] : encrypted_data_buf[1930];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1929] = exp_valid ? exp_out[1929] : encrypted_data_buf[1929];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1928] = exp_valid ? exp_out[1928] : encrypted_data_buf[1928];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1927] = exp_valid ? exp_out[1927] : encrypted_data_buf[1927];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1926] = exp_valid ? exp_out[1926] : encrypted_data_buf[1926];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1925] = exp_valid ? exp_out[1925] : encrypted_data_buf[1925];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1924] = exp_valid ? exp_out[1924] : encrypted_data_buf[1924];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1923] = exp_valid ? exp_out[1923] : encrypted_data_buf[1923];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1922] = exp_valid ? exp_out[1922] : encrypted_data_buf[1922];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1921] = exp_valid ? exp_out[1921] : encrypted_data_buf[1921];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1920] = exp_valid ? exp_out[1920] : encrypted_data_buf[1920];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1919] = exp_valid ? exp_out[1919] : encrypted_data_buf[1919];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1918] = exp_valid ? exp_out[1918] : encrypted_data_buf[1918];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1917] = exp_valid ? exp_out[1917] : encrypted_data_buf[1917];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1916] = exp_valid ? exp_out[1916] : encrypted_data_buf[1916];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1915] = exp_valid ? exp_out[1915] : encrypted_data_buf[1915];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1914] = exp_valid ? exp_out[1914] : encrypted_data_buf[1914];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1913] = exp_valid ? exp_out[1913] : encrypted_data_buf[1913];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1912] = exp_valid ? exp_out[1912] : encrypted_data_buf[1912];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1911] = exp_valid ? exp_out[1911] : encrypted_data_buf[1911];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1910] = exp_valid ? exp_out[1910] : encrypted_data_buf[1910];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1909] = exp_valid ? exp_out[1909] : encrypted_data_buf[1909];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1908] = exp_valid ? exp_out[1908] : encrypted_data_buf[1908];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1907] = exp_valid ? exp_out[1907] : encrypted_data_buf[1907];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1906] = exp_valid ? exp_out[1906] : encrypted_data_buf[1906];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1905] = exp_valid ? exp_out[1905] : encrypted_data_buf[1905];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1904] = exp_valid ? exp_out[1904] : encrypted_data_buf[1904];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1903] = exp_valid ? exp_out[1903] : encrypted_data_buf[1903];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1902] = exp_valid ? exp_out[1902] : encrypted_data_buf[1902];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1901] = exp_valid ? exp_out[1901] : encrypted_data_buf[1901];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1900] = exp_valid ? exp_out[1900] : encrypted_data_buf[1900];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1899] = exp_valid ? exp_out[1899] : encrypted_data_buf[1899];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1898] = exp_valid ? exp_out[1898] : encrypted_data_buf[1898];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1897] = exp_valid ? exp_out[1897] : encrypted_data_buf[1897];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1896] = exp_valid ? exp_out[1896] : encrypted_data_buf[1896];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1895] = exp_valid ? exp_out[1895] : encrypted_data_buf[1895];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1894] = exp_valid ? exp_out[1894] : encrypted_data_buf[1894];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1893] = exp_valid ? exp_out[1893] : encrypted_data_buf[1893];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1892] = exp_valid ? exp_out[1892] : encrypted_data_buf[1892];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1891] = exp_valid ? exp_out[1891] : encrypted_data_buf[1891];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1890] = exp_valid ? exp_out[1890] : encrypted_data_buf[1890];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1889] = exp_valid ? exp_out[1889] : encrypted_data_buf[1889];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1888] = exp_valid ? exp_out[1888] : encrypted_data_buf[1888];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1887] = exp_valid ? exp_out[1887] : encrypted_data_buf[1887];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1886] = exp_valid ? exp_out[1886] : encrypted_data_buf[1886];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1885] = exp_valid ? exp_out[1885] : encrypted_data_buf[1885];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1884] = exp_valid ? exp_out[1884] : encrypted_data_buf[1884];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1883] = exp_valid ? exp_out[1883] : encrypted_data_buf[1883];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1882] = exp_valid ? exp_out[1882] : encrypted_data_buf[1882];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1881] = exp_valid ? exp_out[1881] : encrypted_data_buf[1881];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1880] = exp_valid ? exp_out[1880] : encrypted_data_buf[1880];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1879] = exp_valid ? exp_out[1879] : encrypted_data_buf[1879];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1878] = exp_valid ? exp_out[1878] : encrypted_data_buf[1878];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1877] = exp_valid ? exp_out[1877] : encrypted_data_buf[1877];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1876] = exp_valid ? exp_out[1876] : encrypted_data_buf[1876];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1875] = exp_valid ? exp_out[1875] : encrypted_data_buf[1875];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1874] = exp_valid ? exp_out[1874] : encrypted_data_buf[1874];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1873] = exp_valid ? exp_out[1873] : encrypted_data_buf[1873];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1872] = exp_valid ? exp_out[1872] : encrypted_data_buf[1872];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1871] = exp_valid ? exp_out[1871] : encrypted_data_buf[1871];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1870] = exp_valid ? exp_out[1870] : encrypted_data_buf[1870];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1869] = exp_valid ? exp_out[1869] : encrypted_data_buf[1869];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1868] = exp_valid ? exp_out[1868] : encrypted_data_buf[1868];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1867] = exp_valid ? exp_out[1867] : encrypted_data_buf[1867];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1866] = exp_valid ? exp_out[1866] : encrypted_data_buf[1866];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1865] = exp_valid ? exp_out[1865] : encrypted_data_buf[1865];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1864] = exp_valid ? exp_out[1864] : encrypted_data_buf[1864];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1863] = exp_valid ? exp_out[1863] : encrypted_data_buf[1863];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1862] = exp_valid ? exp_out[1862] : encrypted_data_buf[1862];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1861] = exp_valid ? exp_out[1861] : encrypted_data_buf[1861];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1860] = exp_valid ? exp_out[1860] : encrypted_data_buf[1860];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1859] = exp_valid ? exp_out[1859] : encrypted_data_buf[1859];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1858] = exp_valid ? exp_out[1858] : encrypted_data_buf[1858];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1857] = exp_valid ? exp_out[1857] : encrypted_data_buf[1857];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1856] = exp_valid ? exp_out[1856] : encrypted_data_buf[1856];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1855] = exp_valid ? exp_out[1855] : encrypted_data_buf[1855];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1854] = exp_valid ? exp_out[1854] : encrypted_data_buf[1854];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1853] = exp_valid ? exp_out[1853] : encrypted_data_buf[1853];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1852] = exp_valid ? exp_out[1852] : encrypted_data_buf[1852];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1851] = exp_valid ? exp_out[1851] : encrypted_data_buf[1851];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1850] = exp_valid ? exp_out[1850] : encrypted_data_buf[1850];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1849] = exp_valid ? exp_out[1849] : encrypted_data_buf[1849];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1848] = exp_valid ? exp_out[1848] : encrypted_data_buf[1848];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1847] = exp_valid ? exp_out[1847] : encrypted_data_buf[1847];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1846] = exp_valid ? exp_out[1846] : encrypted_data_buf[1846];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1845] = exp_valid ? exp_out[1845] : encrypted_data_buf[1845];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1844] = exp_valid ? exp_out[1844] : encrypted_data_buf[1844];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1843] = exp_valid ? exp_out[1843] : encrypted_data_buf[1843];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1842] = exp_valid ? exp_out[1842] : encrypted_data_buf[1842];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1841] = exp_valid ? exp_out[1841] : encrypted_data_buf[1841];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1840] = exp_valid ? exp_out[1840] : encrypted_data_buf[1840];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1839] = exp_valid ? exp_out[1839] : encrypted_data_buf[1839];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1838] = exp_valid ? exp_out[1838] : encrypted_data_buf[1838];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1837] = exp_valid ? exp_out[1837] : encrypted_data_buf[1837];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1836] = exp_valid ? exp_out[1836] : encrypted_data_buf[1836];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1835] = exp_valid ? exp_out[1835] : encrypted_data_buf[1835];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1834] = exp_valid ? exp_out[1834] : encrypted_data_buf[1834];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1833] = exp_valid ? exp_out[1833] : encrypted_data_buf[1833];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1832] = exp_valid ? exp_out[1832] : encrypted_data_buf[1832];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1831] = exp_valid ? exp_out[1831] : encrypted_data_buf[1831];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1830] = exp_valid ? exp_out[1830] : encrypted_data_buf[1830];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1829] = exp_valid ? exp_out[1829] : encrypted_data_buf[1829];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1828] = exp_valid ? exp_out[1828] : encrypted_data_buf[1828];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1827] = exp_valid ? exp_out[1827] : encrypted_data_buf[1827];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1826] = exp_valid ? exp_out[1826] : encrypted_data_buf[1826];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1825] = exp_valid ? exp_out[1825] : encrypted_data_buf[1825];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1824] = exp_valid ? exp_out[1824] : encrypted_data_buf[1824];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1823] = exp_valid ? exp_out[1823] : encrypted_data_buf[1823];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1822] = exp_valid ? exp_out[1822] : encrypted_data_buf[1822];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1821] = exp_valid ? exp_out[1821] : encrypted_data_buf[1821];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1820] = exp_valid ? exp_out[1820] : encrypted_data_buf[1820];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1819] = exp_valid ? exp_out[1819] : encrypted_data_buf[1819];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1818] = exp_valid ? exp_out[1818] : encrypted_data_buf[1818];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1817] = exp_valid ? exp_out[1817] : encrypted_data_buf[1817];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1816] = exp_valid ? exp_out[1816] : encrypted_data_buf[1816];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1815] = exp_valid ? exp_out[1815] : encrypted_data_buf[1815];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1814] = exp_valid ? exp_out[1814] : encrypted_data_buf[1814];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1813] = exp_valid ? exp_out[1813] : encrypted_data_buf[1813];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1812] = exp_valid ? exp_out[1812] : encrypted_data_buf[1812];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1811] = exp_valid ? exp_out[1811] : encrypted_data_buf[1811];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1810] = exp_valid ? exp_out[1810] : encrypted_data_buf[1810];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1809] = exp_valid ? exp_out[1809] : encrypted_data_buf[1809];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1808] = exp_valid ? exp_out[1808] : encrypted_data_buf[1808];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1807] = exp_valid ? exp_out[1807] : encrypted_data_buf[1807];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1806] = exp_valid ? exp_out[1806] : encrypted_data_buf[1806];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1805] = exp_valid ? exp_out[1805] : encrypted_data_buf[1805];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1804] = exp_valid ? exp_out[1804] : encrypted_data_buf[1804];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1803] = exp_valid ? exp_out[1803] : encrypted_data_buf[1803];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1802] = exp_valid ? exp_out[1802] : encrypted_data_buf[1802];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1801] = exp_valid ? exp_out[1801] : encrypted_data_buf[1801];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1800] = exp_valid ? exp_out[1800] : encrypted_data_buf[1800];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1799] = exp_valid ? exp_out[1799] : encrypted_data_buf[1799];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1798] = exp_valid ? exp_out[1798] : encrypted_data_buf[1798];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1797] = exp_valid ? exp_out[1797] : encrypted_data_buf[1797];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1796] = exp_valid ? exp_out[1796] : encrypted_data_buf[1796];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1795] = exp_valid ? exp_out[1795] : encrypted_data_buf[1795];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1794] = exp_valid ? exp_out[1794] : encrypted_data_buf[1794];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1793] = exp_valid ? exp_out[1793] : encrypted_data_buf[1793];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1792] = exp_valid ? exp_out[1792] : encrypted_data_buf[1792];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1791] = exp_valid ? exp_out[1791] : encrypted_data_buf[1791];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1790] = exp_valid ? exp_out[1790] : encrypted_data_buf[1790];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1789] = exp_valid ? exp_out[1789] : encrypted_data_buf[1789];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1788] = exp_valid ? exp_out[1788] : encrypted_data_buf[1788];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1787] = exp_valid ? exp_out[1787] : encrypted_data_buf[1787];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1786] = exp_valid ? exp_out[1786] : encrypted_data_buf[1786];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1785] = exp_valid ? exp_out[1785] : encrypted_data_buf[1785];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1784] = exp_valid ? exp_out[1784] : encrypted_data_buf[1784];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1783] = exp_valid ? exp_out[1783] : encrypted_data_buf[1783];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1782] = exp_valid ? exp_out[1782] : encrypted_data_buf[1782];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1781] = exp_valid ? exp_out[1781] : encrypted_data_buf[1781];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1780] = exp_valid ? exp_out[1780] : encrypted_data_buf[1780];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1779] = exp_valid ? exp_out[1779] : encrypted_data_buf[1779];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1778] = exp_valid ? exp_out[1778] : encrypted_data_buf[1778];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1777] = exp_valid ? exp_out[1777] : encrypted_data_buf[1777];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1776] = exp_valid ? exp_out[1776] : encrypted_data_buf[1776];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1775] = exp_valid ? exp_out[1775] : encrypted_data_buf[1775];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1774] = exp_valid ? exp_out[1774] : encrypted_data_buf[1774];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1773] = exp_valid ? exp_out[1773] : encrypted_data_buf[1773];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1772] = exp_valid ? exp_out[1772] : encrypted_data_buf[1772];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1771] = exp_valid ? exp_out[1771] : encrypted_data_buf[1771];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1770] = exp_valid ? exp_out[1770] : encrypted_data_buf[1770];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1769] = exp_valid ? exp_out[1769] : encrypted_data_buf[1769];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1768] = exp_valid ? exp_out[1768] : encrypted_data_buf[1768];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1767] = exp_valid ? exp_out[1767] : encrypted_data_buf[1767];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1766] = exp_valid ? exp_out[1766] : encrypted_data_buf[1766];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1765] = exp_valid ? exp_out[1765] : encrypted_data_buf[1765];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1764] = exp_valid ? exp_out[1764] : encrypted_data_buf[1764];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1763] = exp_valid ? exp_out[1763] : encrypted_data_buf[1763];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1762] = exp_valid ? exp_out[1762] : encrypted_data_buf[1762];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1761] = exp_valid ? exp_out[1761] : encrypted_data_buf[1761];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1760] = exp_valid ? exp_out[1760] : encrypted_data_buf[1760];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1759] = exp_valid ? exp_out[1759] : encrypted_data_buf[1759];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1758] = exp_valid ? exp_out[1758] : encrypted_data_buf[1758];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1757] = exp_valid ? exp_out[1757] : encrypted_data_buf[1757];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1756] = exp_valid ? exp_out[1756] : encrypted_data_buf[1756];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1755] = exp_valid ? exp_out[1755] : encrypted_data_buf[1755];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1754] = exp_valid ? exp_out[1754] : encrypted_data_buf[1754];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1753] = exp_valid ? exp_out[1753] : encrypted_data_buf[1753];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1752] = exp_valid ? exp_out[1752] : encrypted_data_buf[1752];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1751] = exp_valid ? exp_out[1751] : encrypted_data_buf[1751];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1750] = exp_valid ? exp_out[1750] : encrypted_data_buf[1750];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1749] = exp_valid ? exp_out[1749] : encrypted_data_buf[1749];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1748] = exp_valid ? exp_out[1748] : encrypted_data_buf[1748];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1747] = exp_valid ? exp_out[1747] : encrypted_data_buf[1747];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1746] = exp_valid ? exp_out[1746] : encrypted_data_buf[1746];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1745] = exp_valid ? exp_out[1745] : encrypted_data_buf[1745];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1744] = exp_valid ? exp_out[1744] : encrypted_data_buf[1744];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1743] = exp_valid ? exp_out[1743] : encrypted_data_buf[1743];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1742] = exp_valid ? exp_out[1742] : encrypted_data_buf[1742];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1741] = exp_valid ? exp_out[1741] : encrypted_data_buf[1741];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1740] = exp_valid ? exp_out[1740] : encrypted_data_buf[1740];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1739] = exp_valid ? exp_out[1739] : encrypted_data_buf[1739];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1738] = exp_valid ? exp_out[1738] : encrypted_data_buf[1738];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1737] = exp_valid ? exp_out[1737] : encrypted_data_buf[1737];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1736] = exp_valid ? exp_out[1736] : encrypted_data_buf[1736];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1735] = exp_valid ? exp_out[1735] : encrypted_data_buf[1735];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1734] = exp_valid ? exp_out[1734] : encrypted_data_buf[1734];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1733] = exp_valid ? exp_out[1733] : encrypted_data_buf[1733];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1732] = exp_valid ? exp_out[1732] : encrypted_data_buf[1732];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1731] = exp_valid ? exp_out[1731] : encrypted_data_buf[1731];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1730] = exp_valid ? exp_out[1730] : encrypted_data_buf[1730];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1729] = exp_valid ? exp_out[1729] : encrypted_data_buf[1729];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1728] = exp_valid ? exp_out[1728] : encrypted_data_buf[1728];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1727] = exp_valid ? exp_out[1727] : encrypted_data_buf[1727];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1726] = exp_valid ? exp_out[1726] : encrypted_data_buf[1726];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1725] = exp_valid ? exp_out[1725] : encrypted_data_buf[1725];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1724] = exp_valid ? exp_out[1724] : encrypted_data_buf[1724];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1723] = exp_valid ? exp_out[1723] : encrypted_data_buf[1723];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1722] = exp_valid ? exp_out[1722] : encrypted_data_buf[1722];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1721] = exp_valid ? exp_out[1721] : encrypted_data_buf[1721];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1720] = exp_valid ? exp_out[1720] : encrypted_data_buf[1720];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1719] = exp_valid ? exp_out[1719] : encrypted_data_buf[1719];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1718] = exp_valid ? exp_out[1718] : encrypted_data_buf[1718];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1717] = exp_valid ? exp_out[1717] : encrypted_data_buf[1717];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1716] = exp_valid ? exp_out[1716] : encrypted_data_buf[1716];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1715] = exp_valid ? exp_out[1715] : encrypted_data_buf[1715];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1714] = exp_valid ? exp_out[1714] : encrypted_data_buf[1714];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1713] = exp_valid ? exp_out[1713] : encrypted_data_buf[1713];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1712] = exp_valid ? exp_out[1712] : encrypted_data_buf[1712];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1711] = exp_valid ? exp_out[1711] : encrypted_data_buf[1711];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1710] = exp_valid ? exp_out[1710] : encrypted_data_buf[1710];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1709] = exp_valid ? exp_out[1709] : encrypted_data_buf[1709];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1708] = exp_valid ? exp_out[1708] : encrypted_data_buf[1708];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1707] = exp_valid ? exp_out[1707] : encrypted_data_buf[1707];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1706] = exp_valid ? exp_out[1706] : encrypted_data_buf[1706];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1705] = exp_valid ? exp_out[1705] : encrypted_data_buf[1705];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1704] = exp_valid ? exp_out[1704] : encrypted_data_buf[1704];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1703] = exp_valid ? exp_out[1703] : encrypted_data_buf[1703];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1702] = exp_valid ? exp_out[1702] : encrypted_data_buf[1702];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1701] = exp_valid ? exp_out[1701] : encrypted_data_buf[1701];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1700] = exp_valid ? exp_out[1700] : encrypted_data_buf[1700];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1699] = exp_valid ? exp_out[1699] : encrypted_data_buf[1699];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1698] = exp_valid ? exp_out[1698] : encrypted_data_buf[1698];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1697] = exp_valid ? exp_out[1697] : encrypted_data_buf[1697];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1696] = exp_valid ? exp_out[1696] : encrypted_data_buf[1696];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1695] = exp_valid ? exp_out[1695] : encrypted_data_buf[1695];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1694] = exp_valid ? exp_out[1694] : encrypted_data_buf[1694];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1693] = exp_valid ? exp_out[1693] : encrypted_data_buf[1693];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1692] = exp_valid ? exp_out[1692] : encrypted_data_buf[1692];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1691] = exp_valid ? exp_out[1691] : encrypted_data_buf[1691];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1690] = exp_valid ? exp_out[1690] : encrypted_data_buf[1690];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1689] = exp_valid ? exp_out[1689] : encrypted_data_buf[1689];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1688] = exp_valid ? exp_out[1688] : encrypted_data_buf[1688];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1687] = exp_valid ? exp_out[1687] : encrypted_data_buf[1687];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1686] = exp_valid ? exp_out[1686] : encrypted_data_buf[1686];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1685] = exp_valid ? exp_out[1685] : encrypted_data_buf[1685];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1684] = exp_valid ? exp_out[1684] : encrypted_data_buf[1684];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1683] = exp_valid ? exp_out[1683] : encrypted_data_buf[1683];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1682] = exp_valid ? exp_out[1682] : encrypted_data_buf[1682];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1681] = exp_valid ? exp_out[1681] : encrypted_data_buf[1681];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1680] = exp_valid ? exp_out[1680] : encrypted_data_buf[1680];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1679] = exp_valid ? exp_out[1679] : encrypted_data_buf[1679];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1678] = exp_valid ? exp_out[1678] : encrypted_data_buf[1678];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1677] = exp_valid ? exp_out[1677] : encrypted_data_buf[1677];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1676] = exp_valid ? exp_out[1676] : encrypted_data_buf[1676];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1675] = exp_valid ? exp_out[1675] : encrypted_data_buf[1675];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1674] = exp_valid ? exp_out[1674] : encrypted_data_buf[1674];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1673] = exp_valid ? exp_out[1673] : encrypted_data_buf[1673];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1672] = exp_valid ? exp_out[1672] : encrypted_data_buf[1672];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1671] = exp_valid ? exp_out[1671] : encrypted_data_buf[1671];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1670] = exp_valid ? exp_out[1670] : encrypted_data_buf[1670];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1669] = exp_valid ? exp_out[1669] : encrypted_data_buf[1669];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1668] = exp_valid ? exp_out[1668] : encrypted_data_buf[1668];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1667] = exp_valid ? exp_out[1667] : encrypted_data_buf[1667];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1666] = exp_valid ? exp_out[1666] : encrypted_data_buf[1666];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1665] = exp_valid ? exp_out[1665] : encrypted_data_buf[1665];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1664] = exp_valid ? exp_out[1664] : encrypted_data_buf[1664];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1663] = exp_valid ? exp_out[1663] : encrypted_data_buf[1663];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1662] = exp_valid ? exp_out[1662] : encrypted_data_buf[1662];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1661] = exp_valid ? exp_out[1661] : encrypted_data_buf[1661];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1660] = exp_valid ? exp_out[1660] : encrypted_data_buf[1660];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1659] = exp_valid ? exp_out[1659] : encrypted_data_buf[1659];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1658] = exp_valid ? exp_out[1658] : encrypted_data_buf[1658];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1657] = exp_valid ? exp_out[1657] : encrypted_data_buf[1657];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1656] = exp_valid ? exp_out[1656] : encrypted_data_buf[1656];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1655] = exp_valid ? exp_out[1655] : encrypted_data_buf[1655];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1654] = exp_valid ? exp_out[1654] : encrypted_data_buf[1654];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1653] = exp_valid ? exp_out[1653] : encrypted_data_buf[1653];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1652] = exp_valid ? exp_out[1652] : encrypted_data_buf[1652];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1651] = exp_valid ? exp_out[1651] : encrypted_data_buf[1651];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1650] = exp_valid ? exp_out[1650] : encrypted_data_buf[1650];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1649] = exp_valid ? exp_out[1649] : encrypted_data_buf[1649];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1648] = exp_valid ? exp_out[1648] : encrypted_data_buf[1648];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1647] = exp_valid ? exp_out[1647] : encrypted_data_buf[1647];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1646] = exp_valid ? exp_out[1646] : encrypted_data_buf[1646];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1645] = exp_valid ? exp_out[1645] : encrypted_data_buf[1645];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1644] = exp_valid ? exp_out[1644] : encrypted_data_buf[1644];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1643] = exp_valid ? exp_out[1643] : encrypted_data_buf[1643];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1642] = exp_valid ? exp_out[1642] : encrypted_data_buf[1642];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1641] = exp_valid ? exp_out[1641] : encrypted_data_buf[1641];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1640] = exp_valid ? exp_out[1640] : encrypted_data_buf[1640];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1639] = exp_valid ? exp_out[1639] : encrypted_data_buf[1639];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1638] = exp_valid ? exp_out[1638] : encrypted_data_buf[1638];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1637] = exp_valid ? exp_out[1637] : encrypted_data_buf[1637];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1636] = exp_valid ? exp_out[1636] : encrypted_data_buf[1636];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1635] = exp_valid ? exp_out[1635] : encrypted_data_buf[1635];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1634] = exp_valid ? exp_out[1634] : encrypted_data_buf[1634];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1633] = exp_valid ? exp_out[1633] : encrypted_data_buf[1633];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1632] = exp_valid ? exp_out[1632] : encrypted_data_buf[1632];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1631] = exp_valid ? exp_out[1631] : encrypted_data_buf[1631];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1630] = exp_valid ? exp_out[1630] : encrypted_data_buf[1630];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1629] = exp_valid ? exp_out[1629] : encrypted_data_buf[1629];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1628] = exp_valid ? exp_out[1628] : encrypted_data_buf[1628];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1627] = exp_valid ? exp_out[1627] : encrypted_data_buf[1627];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1626] = exp_valid ? exp_out[1626] : encrypted_data_buf[1626];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1625] = exp_valid ? exp_out[1625] : encrypted_data_buf[1625];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1624] = exp_valid ? exp_out[1624] : encrypted_data_buf[1624];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1623] = exp_valid ? exp_out[1623] : encrypted_data_buf[1623];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1622] = exp_valid ? exp_out[1622] : encrypted_data_buf[1622];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1621] = exp_valid ? exp_out[1621] : encrypted_data_buf[1621];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1620] = exp_valid ? exp_out[1620] : encrypted_data_buf[1620];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1619] = exp_valid ? exp_out[1619] : encrypted_data_buf[1619];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1618] = exp_valid ? exp_out[1618] : encrypted_data_buf[1618];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1617] = exp_valid ? exp_out[1617] : encrypted_data_buf[1617];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1616] = exp_valid ? exp_out[1616] : encrypted_data_buf[1616];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1615] = exp_valid ? exp_out[1615] : encrypted_data_buf[1615];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1614] = exp_valid ? exp_out[1614] : encrypted_data_buf[1614];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1613] = exp_valid ? exp_out[1613] : encrypted_data_buf[1613];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1612] = exp_valid ? exp_out[1612] : encrypted_data_buf[1612];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1611] = exp_valid ? exp_out[1611] : encrypted_data_buf[1611];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1610] = exp_valid ? exp_out[1610] : encrypted_data_buf[1610];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1609] = exp_valid ? exp_out[1609] : encrypted_data_buf[1609];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1608] = exp_valid ? exp_out[1608] : encrypted_data_buf[1608];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1607] = exp_valid ? exp_out[1607] : encrypted_data_buf[1607];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1606] = exp_valid ? exp_out[1606] : encrypted_data_buf[1606];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1605] = exp_valid ? exp_out[1605] : encrypted_data_buf[1605];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1604] = exp_valid ? exp_out[1604] : encrypted_data_buf[1604];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1603] = exp_valid ? exp_out[1603] : encrypted_data_buf[1603];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1602] = exp_valid ? exp_out[1602] : encrypted_data_buf[1602];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1601] = exp_valid ? exp_out[1601] : encrypted_data_buf[1601];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1600] = exp_valid ? exp_out[1600] : encrypted_data_buf[1600];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1599] = exp_valid ? exp_out[1599] : encrypted_data_buf[1599];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1598] = exp_valid ? exp_out[1598] : encrypted_data_buf[1598];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1597] = exp_valid ? exp_out[1597] : encrypted_data_buf[1597];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1596] = exp_valid ? exp_out[1596] : encrypted_data_buf[1596];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1595] = exp_valid ? exp_out[1595] : encrypted_data_buf[1595];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1594] = exp_valid ? exp_out[1594] : encrypted_data_buf[1594];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1593] = exp_valid ? exp_out[1593] : encrypted_data_buf[1593];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1592] = exp_valid ? exp_out[1592] : encrypted_data_buf[1592];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1591] = exp_valid ? exp_out[1591] : encrypted_data_buf[1591];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1590] = exp_valid ? exp_out[1590] : encrypted_data_buf[1590];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1589] = exp_valid ? exp_out[1589] : encrypted_data_buf[1589];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1588] = exp_valid ? exp_out[1588] : encrypted_data_buf[1588];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1587] = exp_valid ? exp_out[1587] : encrypted_data_buf[1587];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1586] = exp_valid ? exp_out[1586] : encrypted_data_buf[1586];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1585] = exp_valid ? exp_out[1585] : encrypted_data_buf[1585];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1584] = exp_valid ? exp_out[1584] : encrypted_data_buf[1584];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1583] = exp_valid ? exp_out[1583] : encrypted_data_buf[1583];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1582] = exp_valid ? exp_out[1582] : encrypted_data_buf[1582];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1581] = exp_valid ? exp_out[1581] : encrypted_data_buf[1581];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1580] = exp_valid ? exp_out[1580] : encrypted_data_buf[1580];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1579] = exp_valid ? exp_out[1579] : encrypted_data_buf[1579];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1578] = exp_valid ? exp_out[1578] : encrypted_data_buf[1578];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1577] = exp_valid ? exp_out[1577] : encrypted_data_buf[1577];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1576] = exp_valid ? exp_out[1576] : encrypted_data_buf[1576];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1575] = exp_valid ? exp_out[1575] : encrypted_data_buf[1575];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1574] = exp_valid ? exp_out[1574] : encrypted_data_buf[1574];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1573] = exp_valid ? exp_out[1573] : encrypted_data_buf[1573];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1572] = exp_valid ? exp_out[1572] : encrypted_data_buf[1572];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1571] = exp_valid ? exp_out[1571] : encrypted_data_buf[1571];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1570] = exp_valid ? exp_out[1570] : encrypted_data_buf[1570];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1569] = exp_valid ? exp_out[1569] : encrypted_data_buf[1569];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1568] = exp_valid ? exp_out[1568] : encrypted_data_buf[1568];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1567] = exp_valid ? exp_out[1567] : encrypted_data_buf[1567];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1566] = exp_valid ? exp_out[1566] : encrypted_data_buf[1566];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1565] = exp_valid ? exp_out[1565] : encrypted_data_buf[1565];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1564] = exp_valid ? exp_out[1564] : encrypted_data_buf[1564];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1563] = exp_valid ? exp_out[1563] : encrypted_data_buf[1563];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1562] = exp_valid ? exp_out[1562] : encrypted_data_buf[1562];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1561] = exp_valid ? exp_out[1561] : encrypted_data_buf[1561];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1560] = exp_valid ? exp_out[1560] : encrypted_data_buf[1560];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1559] = exp_valid ? exp_out[1559] : encrypted_data_buf[1559];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1558] = exp_valid ? exp_out[1558] : encrypted_data_buf[1558];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1557] = exp_valid ? exp_out[1557] : encrypted_data_buf[1557];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1556] = exp_valid ? exp_out[1556] : encrypted_data_buf[1556];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1555] = exp_valid ? exp_out[1555] : encrypted_data_buf[1555];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1554] = exp_valid ? exp_out[1554] : encrypted_data_buf[1554];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1553] = exp_valid ? exp_out[1553] : encrypted_data_buf[1553];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1552] = exp_valid ? exp_out[1552] : encrypted_data_buf[1552];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1551] = exp_valid ? exp_out[1551] : encrypted_data_buf[1551];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1550] = exp_valid ? exp_out[1550] : encrypted_data_buf[1550];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1549] = exp_valid ? exp_out[1549] : encrypted_data_buf[1549];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1548] = exp_valid ? exp_out[1548] : encrypted_data_buf[1548];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1547] = exp_valid ? exp_out[1547] : encrypted_data_buf[1547];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1546] = exp_valid ? exp_out[1546] : encrypted_data_buf[1546];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1545] = exp_valid ? exp_out[1545] : encrypted_data_buf[1545];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1544] = exp_valid ? exp_out[1544] : encrypted_data_buf[1544];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1543] = exp_valid ? exp_out[1543] : encrypted_data_buf[1543];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1542] = exp_valid ? exp_out[1542] : encrypted_data_buf[1542];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1541] = exp_valid ? exp_out[1541] : encrypted_data_buf[1541];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1540] = exp_valid ? exp_out[1540] : encrypted_data_buf[1540];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1539] = exp_valid ? exp_out[1539] : encrypted_data_buf[1539];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1538] = exp_valid ? exp_out[1538] : encrypted_data_buf[1538];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1537] = exp_valid ? exp_out[1537] : encrypted_data_buf[1537];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1536] = exp_valid ? exp_out[1536] : encrypted_data_buf[1536];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1535] = exp_valid ? exp_out[1535] : encrypted_data_buf[1535];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1534] = exp_valid ? exp_out[1534] : encrypted_data_buf[1534];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1533] = exp_valid ? exp_out[1533] : encrypted_data_buf[1533];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1532] = exp_valid ? exp_out[1532] : encrypted_data_buf[1532];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1531] = exp_valid ? exp_out[1531] : encrypted_data_buf[1531];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1530] = exp_valid ? exp_out[1530] : encrypted_data_buf[1530];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1529] = exp_valid ? exp_out[1529] : encrypted_data_buf[1529];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1528] = exp_valid ? exp_out[1528] : encrypted_data_buf[1528];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1527] = exp_valid ? exp_out[1527] : encrypted_data_buf[1527];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1526] = exp_valid ? exp_out[1526] : encrypted_data_buf[1526];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1525] = exp_valid ? exp_out[1525] : encrypted_data_buf[1525];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1524] = exp_valid ? exp_out[1524] : encrypted_data_buf[1524];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1523] = exp_valid ? exp_out[1523] : encrypted_data_buf[1523];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1522] = exp_valid ? exp_out[1522] : encrypted_data_buf[1522];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1521] = exp_valid ? exp_out[1521] : encrypted_data_buf[1521];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1520] = exp_valid ? exp_out[1520] : encrypted_data_buf[1520];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1519] = exp_valid ? exp_out[1519] : encrypted_data_buf[1519];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1518] = exp_valid ? exp_out[1518] : encrypted_data_buf[1518];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1517] = exp_valid ? exp_out[1517] : encrypted_data_buf[1517];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1516] = exp_valid ? exp_out[1516] : encrypted_data_buf[1516];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1515] = exp_valid ? exp_out[1515] : encrypted_data_buf[1515];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1514] = exp_valid ? exp_out[1514] : encrypted_data_buf[1514];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1513] = exp_valid ? exp_out[1513] : encrypted_data_buf[1513];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1512] = exp_valid ? exp_out[1512] : encrypted_data_buf[1512];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1511] = exp_valid ? exp_out[1511] : encrypted_data_buf[1511];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1510] = exp_valid ? exp_out[1510] : encrypted_data_buf[1510];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1509] = exp_valid ? exp_out[1509] : encrypted_data_buf[1509];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1508] = exp_valid ? exp_out[1508] : encrypted_data_buf[1508];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1507] = exp_valid ? exp_out[1507] : encrypted_data_buf[1507];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1506] = exp_valid ? exp_out[1506] : encrypted_data_buf[1506];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1505] = exp_valid ? exp_out[1505] : encrypted_data_buf[1505];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1504] = exp_valid ? exp_out[1504] : encrypted_data_buf[1504];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1503] = exp_valid ? exp_out[1503] : encrypted_data_buf[1503];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1502] = exp_valid ? exp_out[1502] : encrypted_data_buf[1502];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1501] = exp_valid ? exp_out[1501] : encrypted_data_buf[1501];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1500] = exp_valid ? exp_out[1500] : encrypted_data_buf[1500];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1499] = exp_valid ? exp_out[1499] : encrypted_data_buf[1499];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1498] = exp_valid ? exp_out[1498] : encrypted_data_buf[1498];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1497] = exp_valid ? exp_out[1497] : encrypted_data_buf[1497];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1496] = exp_valid ? exp_out[1496] : encrypted_data_buf[1496];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1495] = exp_valid ? exp_out[1495] : encrypted_data_buf[1495];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1494] = exp_valid ? exp_out[1494] : encrypted_data_buf[1494];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1493] = exp_valid ? exp_out[1493] : encrypted_data_buf[1493];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1492] = exp_valid ? exp_out[1492] : encrypted_data_buf[1492];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1491] = exp_valid ? exp_out[1491] : encrypted_data_buf[1491];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1490] = exp_valid ? exp_out[1490] : encrypted_data_buf[1490];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1489] = exp_valid ? exp_out[1489] : encrypted_data_buf[1489];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1488] = exp_valid ? exp_out[1488] : encrypted_data_buf[1488];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1487] = exp_valid ? exp_out[1487] : encrypted_data_buf[1487];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1486] = exp_valid ? exp_out[1486] : encrypted_data_buf[1486];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1485] = exp_valid ? exp_out[1485] : encrypted_data_buf[1485];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1484] = exp_valid ? exp_out[1484] : encrypted_data_buf[1484];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1483] = exp_valid ? exp_out[1483] : encrypted_data_buf[1483];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1482] = exp_valid ? exp_out[1482] : encrypted_data_buf[1482];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1481] = exp_valid ? exp_out[1481] : encrypted_data_buf[1481];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1480] = exp_valid ? exp_out[1480] : encrypted_data_buf[1480];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1479] = exp_valid ? exp_out[1479] : encrypted_data_buf[1479];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1478] = exp_valid ? exp_out[1478] : encrypted_data_buf[1478];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1477] = exp_valid ? exp_out[1477] : encrypted_data_buf[1477];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1476] = exp_valid ? exp_out[1476] : encrypted_data_buf[1476];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1475] = exp_valid ? exp_out[1475] : encrypted_data_buf[1475];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1474] = exp_valid ? exp_out[1474] : encrypted_data_buf[1474];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1473] = exp_valid ? exp_out[1473] : encrypted_data_buf[1473];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1472] = exp_valid ? exp_out[1472] : encrypted_data_buf[1472];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1471] = exp_valid ? exp_out[1471] : encrypted_data_buf[1471];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1470] = exp_valid ? exp_out[1470] : encrypted_data_buf[1470];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1469] = exp_valid ? exp_out[1469] : encrypted_data_buf[1469];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1468] = exp_valid ? exp_out[1468] : encrypted_data_buf[1468];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1467] = exp_valid ? exp_out[1467] : encrypted_data_buf[1467];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1466] = exp_valid ? exp_out[1466] : encrypted_data_buf[1466];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1465] = exp_valid ? exp_out[1465] : encrypted_data_buf[1465];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1464] = exp_valid ? exp_out[1464] : encrypted_data_buf[1464];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1463] = exp_valid ? exp_out[1463] : encrypted_data_buf[1463];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1462] = exp_valid ? exp_out[1462] : encrypted_data_buf[1462];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1461] = exp_valid ? exp_out[1461] : encrypted_data_buf[1461];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1460] = exp_valid ? exp_out[1460] : encrypted_data_buf[1460];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1459] = exp_valid ? exp_out[1459] : encrypted_data_buf[1459];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1458] = exp_valid ? exp_out[1458] : encrypted_data_buf[1458];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1457] = exp_valid ? exp_out[1457] : encrypted_data_buf[1457];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1456] = exp_valid ? exp_out[1456] : encrypted_data_buf[1456];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1455] = exp_valid ? exp_out[1455] : encrypted_data_buf[1455];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1454] = exp_valid ? exp_out[1454] : encrypted_data_buf[1454];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1453] = exp_valid ? exp_out[1453] : encrypted_data_buf[1453];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1452] = exp_valid ? exp_out[1452] : encrypted_data_buf[1452];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1451] = exp_valid ? exp_out[1451] : encrypted_data_buf[1451];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1450] = exp_valid ? exp_out[1450] : encrypted_data_buf[1450];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1449] = exp_valid ? exp_out[1449] : encrypted_data_buf[1449];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1448] = exp_valid ? exp_out[1448] : encrypted_data_buf[1448];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1447] = exp_valid ? exp_out[1447] : encrypted_data_buf[1447];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1446] = exp_valid ? exp_out[1446] : encrypted_data_buf[1446];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1445] = exp_valid ? exp_out[1445] : encrypted_data_buf[1445];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1444] = exp_valid ? exp_out[1444] : encrypted_data_buf[1444];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1443] = exp_valid ? exp_out[1443] : encrypted_data_buf[1443];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1442] = exp_valid ? exp_out[1442] : encrypted_data_buf[1442];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1441] = exp_valid ? exp_out[1441] : encrypted_data_buf[1441];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1440] = exp_valid ? exp_out[1440] : encrypted_data_buf[1440];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1439] = exp_valid ? exp_out[1439] : encrypted_data_buf[1439];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1438] = exp_valid ? exp_out[1438] : encrypted_data_buf[1438];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1437] = exp_valid ? exp_out[1437] : encrypted_data_buf[1437];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1436] = exp_valid ? exp_out[1436] : encrypted_data_buf[1436];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1435] = exp_valid ? exp_out[1435] : encrypted_data_buf[1435];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1434] = exp_valid ? exp_out[1434] : encrypted_data_buf[1434];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1433] = exp_valid ? exp_out[1433] : encrypted_data_buf[1433];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1432] = exp_valid ? exp_out[1432] : encrypted_data_buf[1432];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1431] = exp_valid ? exp_out[1431] : encrypted_data_buf[1431];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1430] = exp_valid ? exp_out[1430] : encrypted_data_buf[1430];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1429] = exp_valid ? exp_out[1429] : encrypted_data_buf[1429];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1428] = exp_valid ? exp_out[1428] : encrypted_data_buf[1428];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1427] = exp_valid ? exp_out[1427] : encrypted_data_buf[1427];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1426] = exp_valid ? exp_out[1426] : encrypted_data_buf[1426];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1425] = exp_valid ? exp_out[1425] : encrypted_data_buf[1425];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1424] = exp_valid ? exp_out[1424] : encrypted_data_buf[1424];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1423] = exp_valid ? exp_out[1423] : encrypted_data_buf[1423];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1422] = exp_valid ? exp_out[1422] : encrypted_data_buf[1422];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1421] = exp_valid ? exp_out[1421] : encrypted_data_buf[1421];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1420] = exp_valid ? exp_out[1420] : encrypted_data_buf[1420];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1419] = exp_valid ? exp_out[1419] : encrypted_data_buf[1419];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1418] = exp_valid ? exp_out[1418] : encrypted_data_buf[1418];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1417] = exp_valid ? exp_out[1417] : encrypted_data_buf[1417];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1416] = exp_valid ? exp_out[1416] : encrypted_data_buf[1416];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1415] = exp_valid ? exp_out[1415] : encrypted_data_buf[1415];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1414] = exp_valid ? exp_out[1414] : encrypted_data_buf[1414];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1413] = exp_valid ? exp_out[1413] : encrypted_data_buf[1413];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1412] = exp_valid ? exp_out[1412] : encrypted_data_buf[1412];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1411] = exp_valid ? exp_out[1411] : encrypted_data_buf[1411];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1410] = exp_valid ? exp_out[1410] : encrypted_data_buf[1410];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1409] = exp_valid ? exp_out[1409] : encrypted_data_buf[1409];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1408] = exp_valid ? exp_out[1408] : encrypted_data_buf[1408];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1407] = exp_valid ? exp_out[1407] : encrypted_data_buf[1407];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1406] = exp_valid ? exp_out[1406] : encrypted_data_buf[1406];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1405] = exp_valid ? exp_out[1405] : encrypted_data_buf[1405];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1404] = exp_valid ? exp_out[1404] : encrypted_data_buf[1404];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1403] = exp_valid ? exp_out[1403] : encrypted_data_buf[1403];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1402] = exp_valid ? exp_out[1402] : encrypted_data_buf[1402];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1401] = exp_valid ? exp_out[1401] : encrypted_data_buf[1401];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1400] = exp_valid ? exp_out[1400] : encrypted_data_buf[1400];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1399] = exp_valid ? exp_out[1399] : encrypted_data_buf[1399];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1398] = exp_valid ? exp_out[1398] : encrypted_data_buf[1398];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1397] = exp_valid ? exp_out[1397] : encrypted_data_buf[1397];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1396] = exp_valid ? exp_out[1396] : encrypted_data_buf[1396];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1395] = exp_valid ? exp_out[1395] : encrypted_data_buf[1395];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1394] = exp_valid ? exp_out[1394] : encrypted_data_buf[1394];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1393] = exp_valid ? exp_out[1393] : encrypted_data_buf[1393];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1392] = exp_valid ? exp_out[1392] : encrypted_data_buf[1392];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1391] = exp_valid ? exp_out[1391] : encrypted_data_buf[1391];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1390] = exp_valid ? exp_out[1390] : encrypted_data_buf[1390];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1389] = exp_valid ? exp_out[1389] : encrypted_data_buf[1389];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1388] = exp_valid ? exp_out[1388] : encrypted_data_buf[1388];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1387] = exp_valid ? exp_out[1387] : encrypted_data_buf[1387];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1386] = exp_valid ? exp_out[1386] : encrypted_data_buf[1386];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1385] = exp_valid ? exp_out[1385] : encrypted_data_buf[1385];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1384] = exp_valid ? exp_out[1384] : encrypted_data_buf[1384];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1383] = exp_valid ? exp_out[1383] : encrypted_data_buf[1383];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1382] = exp_valid ? exp_out[1382] : encrypted_data_buf[1382];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1381] = exp_valid ? exp_out[1381] : encrypted_data_buf[1381];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1380] = exp_valid ? exp_out[1380] : encrypted_data_buf[1380];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1379] = exp_valid ? exp_out[1379] : encrypted_data_buf[1379];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1378] = exp_valid ? exp_out[1378] : encrypted_data_buf[1378];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1377] = exp_valid ? exp_out[1377] : encrypted_data_buf[1377];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1376] = exp_valid ? exp_out[1376] : encrypted_data_buf[1376];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1375] = exp_valid ? exp_out[1375] : encrypted_data_buf[1375];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1374] = exp_valid ? exp_out[1374] : encrypted_data_buf[1374];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1373] = exp_valid ? exp_out[1373] : encrypted_data_buf[1373];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1372] = exp_valid ? exp_out[1372] : encrypted_data_buf[1372];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1371] = exp_valid ? exp_out[1371] : encrypted_data_buf[1371];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1370] = exp_valid ? exp_out[1370] : encrypted_data_buf[1370];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1369] = exp_valid ? exp_out[1369] : encrypted_data_buf[1369];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1368] = exp_valid ? exp_out[1368] : encrypted_data_buf[1368];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1367] = exp_valid ? exp_out[1367] : encrypted_data_buf[1367];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1366] = exp_valid ? exp_out[1366] : encrypted_data_buf[1366];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1365] = exp_valid ? exp_out[1365] : encrypted_data_buf[1365];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1364] = exp_valid ? exp_out[1364] : encrypted_data_buf[1364];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1363] = exp_valid ? exp_out[1363] : encrypted_data_buf[1363];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1362] = exp_valid ? exp_out[1362] : encrypted_data_buf[1362];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1361] = exp_valid ? exp_out[1361] : encrypted_data_buf[1361];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1360] = exp_valid ? exp_out[1360] : encrypted_data_buf[1360];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1359] = exp_valid ? exp_out[1359] : encrypted_data_buf[1359];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1358] = exp_valid ? exp_out[1358] : encrypted_data_buf[1358];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1357] = exp_valid ? exp_out[1357] : encrypted_data_buf[1357];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1356] = exp_valid ? exp_out[1356] : encrypted_data_buf[1356];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1355] = exp_valid ? exp_out[1355] : encrypted_data_buf[1355];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1354] = exp_valid ? exp_out[1354] : encrypted_data_buf[1354];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1353] = exp_valid ? exp_out[1353] : encrypted_data_buf[1353];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1352] = exp_valid ? exp_out[1352] : encrypted_data_buf[1352];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1351] = exp_valid ? exp_out[1351] : encrypted_data_buf[1351];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1350] = exp_valid ? exp_out[1350] : encrypted_data_buf[1350];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1349] = exp_valid ? exp_out[1349] : encrypted_data_buf[1349];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1348] = exp_valid ? exp_out[1348] : encrypted_data_buf[1348];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1347] = exp_valid ? exp_out[1347] : encrypted_data_buf[1347];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1346] = exp_valid ? exp_out[1346] : encrypted_data_buf[1346];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1345] = exp_valid ? exp_out[1345] : encrypted_data_buf[1345];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1344] = exp_valid ? exp_out[1344] : encrypted_data_buf[1344];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1343] = exp_valid ? exp_out[1343] : encrypted_data_buf[1343];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1342] = exp_valid ? exp_out[1342] : encrypted_data_buf[1342];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1341] = exp_valid ? exp_out[1341] : encrypted_data_buf[1341];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1340] = exp_valid ? exp_out[1340] : encrypted_data_buf[1340];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1339] = exp_valid ? exp_out[1339] : encrypted_data_buf[1339];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1338] = exp_valid ? exp_out[1338] : encrypted_data_buf[1338];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1337] = exp_valid ? exp_out[1337] : encrypted_data_buf[1337];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1336] = exp_valid ? exp_out[1336] : encrypted_data_buf[1336];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1335] = exp_valid ? exp_out[1335] : encrypted_data_buf[1335];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1334] = exp_valid ? exp_out[1334] : encrypted_data_buf[1334];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1333] = exp_valid ? exp_out[1333] : encrypted_data_buf[1333];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1332] = exp_valid ? exp_out[1332] : encrypted_data_buf[1332];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1331] = exp_valid ? exp_out[1331] : encrypted_data_buf[1331];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1330] = exp_valid ? exp_out[1330] : encrypted_data_buf[1330];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1329] = exp_valid ? exp_out[1329] : encrypted_data_buf[1329];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1328] = exp_valid ? exp_out[1328] : encrypted_data_buf[1328];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1327] = exp_valid ? exp_out[1327] : encrypted_data_buf[1327];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1326] = exp_valid ? exp_out[1326] : encrypted_data_buf[1326];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1325] = exp_valid ? exp_out[1325] : encrypted_data_buf[1325];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1324] = exp_valid ? exp_out[1324] : encrypted_data_buf[1324];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1323] = exp_valid ? exp_out[1323] : encrypted_data_buf[1323];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1322] = exp_valid ? exp_out[1322] : encrypted_data_buf[1322];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1321] = exp_valid ? exp_out[1321] : encrypted_data_buf[1321];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1320] = exp_valid ? exp_out[1320] : encrypted_data_buf[1320];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1319] = exp_valid ? exp_out[1319] : encrypted_data_buf[1319];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1318] = exp_valid ? exp_out[1318] : encrypted_data_buf[1318];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1317] = exp_valid ? exp_out[1317] : encrypted_data_buf[1317];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1316] = exp_valid ? exp_out[1316] : encrypted_data_buf[1316];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1315] = exp_valid ? exp_out[1315] : encrypted_data_buf[1315];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1314] = exp_valid ? exp_out[1314] : encrypted_data_buf[1314];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1313] = exp_valid ? exp_out[1313] : encrypted_data_buf[1313];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1312] = exp_valid ? exp_out[1312] : encrypted_data_buf[1312];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1311] = exp_valid ? exp_out[1311] : encrypted_data_buf[1311];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1310] = exp_valid ? exp_out[1310] : encrypted_data_buf[1310];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1309] = exp_valid ? exp_out[1309] : encrypted_data_buf[1309];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1308] = exp_valid ? exp_out[1308] : encrypted_data_buf[1308];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1307] = exp_valid ? exp_out[1307] : encrypted_data_buf[1307];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1306] = exp_valid ? exp_out[1306] : encrypted_data_buf[1306];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1305] = exp_valid ? exp_out[1305] : encrypted_data_buf[1305];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1304] = exp_valid ? exp_out[1304] : encrypted_data_buf[1304];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1303] = exp_valid ? exp_out[1303] : encrypted_data_buf[1303];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1302] = exp_valid ? exp_out[1302] : encrypted_data_buf[1302];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1301] = exp_valid ? exp_out[1301] : encrypted_data_buf[1301];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1300] = exp_valid ? exp_out[1300] : encrypted_data_buf[1300];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1299] = exp_valid ? exp_out[1299] : encrypted_data_buf[1299];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1298] = exp_valid ? exp_out[1298] : encrypted_data_buf[1298];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1297] = exp_valid ? exp_out[1297] : encrypted_data_buf[1297];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1296] = exp_valid ? exp_out[1296] : encrypted_data_buf[1296];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1295] = exp_valid ? exp_out[1295] : encrypted_data_buf[1295];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1294] = exp_valid ? exp_out[1294] : encrypted_data_buf[1294];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1293] = exp_valid ? exp_out[1293] : encrypted_data_buf[1293];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1292] = exp_valid ? exp_out[1292] : encrypted_data_buf[1292];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1291] = exp_valid ? exp_out[1291] : encrypted_data_buf[1291];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1290] = exp_valid ? exp_out[1290] : encrypted_data_buf[1290];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1289] = exp_valid ? exp_out[1289] : encrypted_data_buf[1289];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1288] = exp_valid ? exp_out[1288] : encrypted_data_buf[1288];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1287] = exp_valid ? exp_out[1287] : encrypted_data_buf[1287];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1286] = exp_valid ? exp_out[1286] : encrypted_data_buf[1286];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1285] = exp_valid ? exp_out[1285] : encrypted_data_buf[1285];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1284] = exp_valid ? exp_out[1284] : encrypted_data_buf[1284];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1283] = exp_valid ? exp_out[1283] : encrypted_data_buf[1283];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1282] = exp_valid ? exp_out[1282] : encrypted_data_buf[1282];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1281] = exp_valid ? exp_out[1281] : encrypted_data_buf[1281];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1280] = exp_valid ? exp_out[1280] : encrypted_data_buf[1280];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1279] = exp_valid ? exp_out[1279] : encrypted_data_buf[1279];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1278] = exp_valid ? exp_out[1278] : encrypted_data_buf[1278];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1277] = exp_valid ? exp_out[1277] : encrypted_data_buf[1277];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1276] = exp_valid ? exp_out[1276] : encrypted_data_buf[1276];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1275] = exp_valid ? exp_out[1275] : encrypted_data_buf[1275];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1274] = exp_valid ? exp_out[1274] : encrypted_data_buf[1274];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1273] = exp_valid ? exp_out[1273] : encrypted_data_buf[1273];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1272] = exp_valid ? exp_out[1272] : encrypted_data_buf[1272];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1271] = exp_valid ? exp_out[1271] : encrypted_data_buf[1271];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1270] = exp_valid ? exp_out[1270] : encrypted_data_buf[1270];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1269] = exp_valid ? exp_out[1269] : encrypted_data_buf[1269];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1268] = exp_valid ? exp_out[1268] : encrypted_data_buf[1268];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1267] = exp_valid ? exp_out[1267] : encrypted_data_buf[1267];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1266] = exp_valid ? exp_out[1266] : encrypted_data_buf[1266];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1265] = exp_valid ? exp_out[1265] : encrypted_data_buf[1265];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1264] = exp_valid ? exp_out[1264] : encrypted_data_buf[1264];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1263] = exp_valid ? exp_out[1263] : encrypted_data_buf[1263];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1262] = exp_valid ? exp_out[1262] : encrypted_data_buf[1262];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1261] = exp_valid ? exp_out[1261] : encrypted_data_buf[1261];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1260] = exp_valid ? exp_out[1260] : encrypted_data_buf[1260];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1259] = exp_valid ? exp_out[1259] : encrypted_data_buf[1259];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1258] = exp_valid ? exp_out[1258] : encrypted_data_buf[1258];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1257] = exp_valid ? exp_out[1257] : encrypted_data_buf[1257];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1256] = exp_valid ? exp_out[1256] : encrypted_data_buf[1256];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1255] = exp_valid ? exp_out[1255] : encrypted_data_buf[1255];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1254] = exp_valid ? exp_out[1254] : encrypted_data_buf[1254];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1253] = exp_valid ? exp_out[1253] : encrypted_data_buf[1253];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1252] = exp_valid ? exp_out[1252] : encrypted_data_buf[1252];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1251] = exp_valid ? exp_out[1251] : encrypted_data_buf[1251];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1250] = exp_valid ? exp_out[1250] : encrypted_data_buf[1250];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1249] = exp_valid ? exp_out[1249] : encrypted_data_buf[1249];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1248] = exp_valid ? exp_out[1248] : encrypted_data_buf[1248];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1247] = exp_valid ? exp_out[1247] : encrypted_data_buf[1247];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1246] = exp_valid ? exp_out[1246] : encrypted_data_buf[1246];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1245] = exp_valid ? exp_out[1245] : encrypted_data_buf[1245];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1244] = exp_valid ? exp_out[1244] : encrypted_data_buf[1244];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1243] = exp_valid ? exp_out[1243] : encrypted_data_buf[1243];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1242] = exp_valid ? exp_out[1242] : encrypted_data_buf[1242];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1241] = exp_valid ? exp_out[1241] : encrypted_data_buf[1241];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1240] = exp_valid ? exp_out[1240] : encrypted_data_buf[1240];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1239] = exp_valid ? exp_out[1239] : encrypted_data_buf[1239];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1238] = exp_valid ? exp_out[1238] : encrypted_data_buf[1238];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1237] = exp_valid ? exp_out[1237] : encrypted_data_buf[1237];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1236] = exp_valid ? exp_out[1236] : encrypted_data_buf[1236];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1235] = exp_valid ? exp_out[1235] : encrypted_data_buf[1235];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1234] = exp_valid ? exp_out[1234] : encrypted_data_buf[1234];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1233] = exp_valid ? exp_out[1233] : encrypted_data_buf[1233];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1232] = exp_valid ? exp_out[1232] : encrypted_data_buf[1232];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1231] = exp_valid ? exp_out[1231] : encrypted_data_buf[1231];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1230] = exp_valid ? exp_out[1230] : encrypted_data_buf[1230];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1229] = exp_valid ? exp_out[1229] : encrypted_data_buf[1229];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1228] = exp_valid ? exp_out[1228] : encrypted_data_buf[1228];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1227] = exp_valid ? exp_out[1227] : encrypted_data_buf[1227];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1226] = exp_valid ? exp_out[1226] : encrypted_data_buf[1226];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1225] = exp_valid ? exp_out[1225] : encrypted_data_buf[1225];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1224] = exp_valid ? exp_out[1224] : encrypted_data_buf[1224];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1223] = exp_valid ? exp_out[1223] : encrypted_data_buf[1223];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1222] = exp_valid ? exp_out[1222] : encrypted_data_buf[1222];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1221] = exp_valid ? exp_out[1221] : encrypted_data_buf[1221];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1220] = exp_valid ? exp_out[1220] : encrypted_data_buf[1220];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1219] = exp_valid ? exp_out[1219] : encrypted_data_buf[1219];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1218] = exp_valid ? exp_out[1218] : encrypted_data_buf[1218];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1217] = exp_valid ? exp_out[1217] : encrypted_data_buf[1217];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1216] = exp_valid ? exp_out[1216] : encrypted_data_buf[1216];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1215] = exp_valid ? exp_out[1215] : encrypted_data_buf[1215];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1214] = exp_valid ? exp_out[1214] : encrypted_data_buf[1214];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1213] = exp_valid ? exp_out[1213] : encrypted_data_buf[1213];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1212] = exp_valid ? exp_out[1212] : encrypted_data_buf[1212];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1211] = exp_valid ? exp_out[1211] : encrypted_data_buf[1211];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1210] = exp_valid ? exp_out[1210] : encrypted_data_buf[1210];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1209] = exp_valid ? exp_out[1209] : encrypted_data_buf[1209];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1208] = exp_valid ? exp_out[1208] : encrypted_data_buf[1208];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1207] = exp_valid ? exp_out[1207] : encrypted_data_buf[1207];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1206] = exp_valid ? exp_out[1206] : encrypted_data_buf[1206];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1205] = exp_valid ? exp_out[1205] : encrypted_data_buf[1205];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1204] = exp_valid ? exp_out[1204] : encrypted_data_buf[1204];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1203] = exp_valid ? exp_out[1203] : encrypted_data_buf[1203];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1202] = exp_valid ? exp_out[1202] : encrypted_data_buf[1202];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1201] = exp_valid ? exp_out[1201] : encrypted_data_buf[1201];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1200] = exp_valid ? exp_out[1200] : encrypted_data_buf[1200];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1199] = exp_valid ? exp_out[1199] : encrypted_data_buf[1199];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1198] = exp_valid ? exp_out[1198] : encrypted_data_buf[1198];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1197] = exp_valid ? exp_out[1197] : encrypted_data_buf[1197];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1196] = exp_valid ? exp_out[1196] : encrypted_data_buf[1196];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1195] = exp_valid ? exp_out[1195] : encrypted_data_buf[1195];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1194] = exp_valid ? exp_out[1194] : encrypted_data_buf[1194];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1193] = exp_valid ? exp_out[1193] : encrypted_data_buf[1193];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1192] = exp_valid ? exp_out[1192] : encrypted_data_buf[1192];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1191] = exp_valid ? exp_out[1191] : encrypted_data_buf[1191];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1190] = exp_valid ? exp_out[1190] : encrypted_data_buf[1190];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1189] = exp_valid ? exp_out[1189] : encrypted_data_buf[1189];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1188] = exp_valid ? exp_out[1188] : encrypted_data_buf[1188];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1187] = exp_valid ? exp_out[1187] : encrypted_data_buf[1187];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1186] = exp_valid ? exp_out[1186] : encrypted_data_buf[1186];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1185] = exp_valid ? exp_out[1185] : encrypted_data_buf[1185];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1184] = exp_valid ? exp_out[1184] : encrypted_data_buf[1184];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1183] = exp_valid ? exp_out[1183] : encrypted_data_buf[1183];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1182] = exp_valid ? exp_out[1182] : encrypted_data_buf[1182];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1181] = exp_valid ? exp_out[1181] : encrypted_data_buf[1181];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1180] = exp_valid ? exp_out[1180] : encrypted_data_buf[1180];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1179] = exp_valid ? exp_out[1179] : encrypted_data_buf[1179];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1178] = exp_valid ? exp_out[1178] : encrypted_data_buf[1178];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1177] = exp_valid ? exp_out[1177] : encrypted_data_buf[1177];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1176] = exp_valid ? exp_out[1176] : encrypted_data_buf[1176];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1175] = exp_valid ? exp_out[1175] : encrypted_data_buf[1175];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1174] = exp_valid ? exp_out[1174] : encrypted_data_buf[1174];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1173] = exp_valid ? exp_out[1173] : encrypted_data_buf[1173];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1172] = exp_valid ? exp_out[1172] : encrypted_data_buf[1172];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1171] = exp_valid ? exp_out[1171] : encrypted_data_buf[1171];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1170] = exp_valid ? exp_out[1170] : encrypted_data_buf[1170];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1169] = exp_valid ? exp_out[1169] : encrypted_data_buf[1169];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1168] = exp_valid ? exp_out[1168] : encrypted_data_buf[1168];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1167] = exp_valid ? exp_out[1167] : encrypted_data_buf[1167];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1166] = exp_valid ? exp_out[1166] : encrypted_data_buf[1166];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1165] = exp_valid ? exp_out[1165] : encrypted_data_buf[1165];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1164] = exp_valid ? exp_out[1164] : encrypted_data_buf[1164];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1163] = exp_valid ? exp_out[1163] : encrypted_data_buf[1163];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1162] = exp_valid ? exp_out[1162] : encrypted_data_buf[1162];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1161] = exp_valid ? exp_out[1161] : encrypted_data_buf[1161];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1160] = exp_valid ? exp_out[1160] : encrypted_data_buf[1160];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1159] = exp_valid ? exp_out[1159] : encrypted_data_buf[1159];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1158] = exp_valid ? exp_out[1158] : encrypted_data_buf[1158];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1157] = exp_valid ? exp_out[1157] : encrypted_data_buf[1157];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1156] = exp_valid ? exp_out[1156] : encrypted_data_buf[1156];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1155] = exp_valid ? exp_out[1155] : encrypted_data_buf[1155];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1154] = exp_valid ? exp_out[1154] : encrypted_data_buf[1154];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1153] = exp_valid ? exp_out[1153] : encrypted_data_buf[1153];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1152] = exp_valid ? exp_out[1152] : encrypted_data_buf[1152];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1151] = exp_valid ? exp_out[1151] : encrypted_data_buf[1151];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1150] = exp_valid ? exp_out[1150] : encrypted_data_buf[1150];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1149] = exp_valid ? exp_out[1149] : encrypted_data_buf[1149];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1148] = exp_valid ? exp_out[1148] : encrypted_data_buf[1148];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1147] = exp_valid ? exp_out[1147] : encrypted_data_buf[1147];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1146] = exp_valid ? exp_out[1146] : encrypted_data_buf[1146];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1145] = exp_valid ? exp_out[1145] : encrypted_data_buf[1145];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1144] = exp_valid ? exp_out[1144] : encrypted_data_buf[1144];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1143] = exp_valid ? exp_out[1143] : encrypted_data_buf[1143];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1142] = exp_valid ? exp_out[1142] : encrypted_data_buf[1142];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1141] = exp_valid ? exp_out[1141] : encrypted_data_buf[1141];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1140] = exp_valid ? exp_out[1140] : encrypted_data_buf[1140];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1139] = exp_valid ? exp_out[1139] : encrypted_data_buf[1139];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1138] = exp_valid ? exp_out[1138] : encrypted_data_buf[1138];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1137] = exp_valid ? exp_out[1137] : encrypted_data_buf[1137];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1136] = exp_valid ? exp_out[1136] : encrypted_data_buf[1136];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1135] = exp_valid ? exp_out[1135] : encrypted_data_buf[1135];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1134] = exp_valid ? exp_out[1134] : encrypted_data_buf[1134];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1133] = exp_valid ? exp_out[1133] : encrypted_data_buf[1133];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1132] = exp_valid ? exp_out[1132] : encrypted_data_buf[1132];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1131] = exp_valid ? exp_out[1131] : encrypted_data_buf[1131];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1130] = exp_valid ? exp_out[1130] : encrypted_data_buf[1130];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1129] = exp_valid ? exp_out[1129] : encrypted_data_buf[1129];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1128] = exp_valid ? exp_out[1128] : encrypted_data_buf[1128];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1127] = exp_valid ? exp_out[1127] : encrypted_data_buf[1127];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1126] = exp_valid ? exp_out[1126] : encrypted_data_buf[1126];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1125] = exp_valid ? exp_out[1125] : encrypted_data_buf[1125];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1124] = exp_valid ? exp_out[1124] : encrypted_data_buf[1124];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1123] = exp_valid ? exp_out[1123] : encrypted_data_buf[1123];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1122] = exp_valid ? exp_out[1122] : encrypted_data_buf[1122];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1121] = exp_valid ? exp_out[1121] : encrypted_data_buf[1121];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1120] = exp_valid ? exp_out[1120] : encrypted_data_buf[1120];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1119] = exp_valid ? exp_out[1119] : encrypted_data_buf[1119];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1118] = exp_valid ? exp_out[1118] : encrypted_data_buf[1118];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1117] = exp_valid ? exp_out[1117] : encrypted_data_buf[1117];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1116] = exp_valid ? exp_out[1116] : encrypted_data_buf[1116];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1115] = exp_valid ? exp_out[1115] : encrypted_data_buf[1115];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1114] = exp_valid ? exp_out[1114] : encrypted_data_buf[1114];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1113] = exp_valid ? exp_out[1113] : encrypted_data_buf[1113];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1112] = exp_valid ? exp_out[1112] : encrypted_data_buf[1112];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1111] = exp_valid ? exp_out[1111] : encrypted_data_buf[1111];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1110] = exp_valid ? exp_out[1110] : encrypted_data_buf[1110];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1109] = exp_valid ? exp_out[1109] : encrypted_data_buf[1109];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1108] = exp_valid ? exp_out[1108] : encrypted_data_buf[1108];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1107] = exp_valid ? exp_out[1107] : encrypted_data_buf[1107];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1106] = exp_valid ? exp_out[1106] : encrypted_data_buf[1106];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1105] = exp_valid ? exp_out[1105] : encrypted_data_buf[1105];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1104] = exp_valid ? exp_out[1104] : encrypted_data_buf[1104];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1103] = exp_valid ? exp_out[1103] : encrypted_data_buf[1103];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1102] = exp_valid ? exp_out[1102] : encrypted_data_buf[1102];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1101] = exp_valid ? exp_out[1101] : encrypted_data_buf[1101];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1100] = exp_valid ? exp_out[1100] : encrypted_data_buf[1100];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1099] = exp_valid ? exp_out[1099] : encrypted_data_buf[1099];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1098] = exp_valid ? exp_out[1098] : encrypted_data_buf[1098];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1097] = exp_valid ? exp_out[1097] : encrypted_data_buf[1097];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1096] = exp_valid ? exp_out[1096] : encrypted_data_buf[1096];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1095] = exp_valid ? exp_out[1095] : encrypted_data_buf[1095];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1094] = exp_valid ? exp_out[1094] : encrypted_data_buf[1094];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1093] = exp_valid ? exp_out[1093] : encrypted_data_buf[1093];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1092] = exp_valid ? exp_out[1092] : encrypted_data_buf[1092];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1091] = exp_valid ? exp_out[1091] : encrypted_data_buf[1091];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1090] = exp_valid ? exp_out[1090] : encrypted_data_buf[1090];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1089] = exp_valid ? exp_out[1089] : encrypted_data_buf[1089];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1088] = exp_valid ? exp_out[1088] : encrypted_data_buf[1088];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1087] = exp_valid ? exp_out[1087] : encrypted_data_buf[1087];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1086] = exp_valid ? exp_out[1086] : encrypted_data_buf[1086];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1085] = exp_valid ? exp_out[1085] : encrypted_data_buf[1085];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1084] = exp_valid ? exp_out[1084] : encrypted_data_buf[1084];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1083] = exp_valid ? exp_out[1083] : encrypted_data_buf[1083];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1082] = exp_valid ? exp_out[1082] : encrypted_data_buf[1082];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1081] = exp_valid ? exp_out[1081] : encrypted_data_buf[1081];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1080] = exp_valid ? exp_out[1080] : encrypted_data_buf[1080];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1079] = exp_valid ? exp_out[1079] : encrypted_data_buf[1079];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1078] = exp_valid ? exp_out[1078] : encrypted_data_buf[1078];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1077] = exp_valid ? exp_out[1077] : encrypted_data_buf[1077];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1076] = exp_valid ? exp_out[1076] : encrypted_data_buf[1076];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1075] = exp_valid ? exp_out[1075] : encrypted_data_buf[1075];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1074] = exp_valid ? exp_out[1074] : encrypted_data_buf[1074];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1073] = exp_valid ? exp_out[1073] : encrypted_data_buf[1073];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1072] = exp_valid ? exp_out[1072] : encrypted_data_buf[1072];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1071] = exp_valid ? exp_out[1071] : encrypted_data_buf[1071];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1070] = exp_valid ? exp_out[1070] : encrypted_data_buf[1070];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1069] = exp_valid ? exp_out[1069] : encrypted_data_buf[1069];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1068] = exp_valid ? exp_out[1068] : encrypted_data_buf[1068];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1067] = exp_valid ? exp_out[1067] : encrypted_data_buf[1067];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1066] = exp_valid ? exp_out[1066] : encrypted_data_buf[1066];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1065] = exp_valid ? exp_out[1065] : encrypted_data_buf[1065];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1064] = exp_valid ? exp_out[1064] : encrypted_data_buf[1064];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1063] = exp_valid ? exp_out[1063] : encrypted_data_buf[1063];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1062] = exp_valid ? exp_out[1062] : encrypted_data_buf[1062];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1061] = exp_valid ? exp_out[1061] : encrypted_data_buf[1061];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1060] = exp_valid ? exp_out[1060] : encrypted_data_buf[1060];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1059] = exp_valid ? exp_out[1059] : encrypted_data_buf[1059];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1058] = exp_valid ? exp_out[1058] : encrypted_data_buf[1058];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1057] = exp_valid ? exp_out[1057] : encrypted_data_buf[1057];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1056] = exp_valid ? exp_out[1056] : encrypted_data_buf[1056];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1055] = exp_valid ? exp_out[1055] : encrypted_data_buf[1055];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1054] = exp_valid ? exp_out[1054] : encrypted_data_buf[1054];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1053] = exp_valid ? exp_out[1053] : encrypted_data_buf[1053];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1052] = exp_valid ? exp_out[1052] : encrypted_data_buf[1052];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1051] = exp_valid ? exp_out[1051] : encrypted_data_buf[1051];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1050] = exp_valid ? exp_out[1050] : encrypted_data_buf[1050];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1049] = exp_valid ? exp_out[1049] : encrypted_data_buf[1049];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1048] = exp_valid ? exp_out[1048] : encrypted_data_buf[1048];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1047] = exp_valid ? exp_out[1047] : encrypted_data_buf[1047];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1046] = exp_valid ? exp_out[1046] : encrypted_data_buf[1046];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1045] = exp_valid ? exp_out[1045] : encrypted_data_buf[1045];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1044] = exp_valid ? exp_out[1044] : encrypted_data_buf[1044];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1043] = exp_valid ? exp_out[1043] : encrypted_data_buf[1043];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1042] = exp_valid ? exp_out[1042] : encrypted_data_buf[1042];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1041] = exp_valid ? exp_out[1041] : encrypted_data_buf[1041];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1040] = exp_valid ? exp_out[1040] : encrypted_data_buf[1040];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1039] = exp_valid ? exp_out[1039] : encrypted_data_buf[1039];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1038] = exp_valid ? exp_out[1038] : encrypted_data_buf[1038];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1037] = exp_valid ? exp_out[1037] : encrypted_data_buf[1037];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1036] = exp_valid ? exp_out[1036] : encrypted_data_buf[1036];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1035] = exp_valid ? exp_out[1035] : encrypted_data_buf[1035];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1034] = exp_valid ? exp_out[1034] : encrypted_data_buf[1034];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1033] = exp_valid ? exp_out[1033] : encrypted_data_buf[1033];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1032] = exp_valid ? exp_out[1032] : encrypted_data_buf[1032];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1031] = exp_valid ? exp_out[1031] : encrypted_data_buf[1031];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1030] = exp_valid ? exp_out[1030] : encrypted_data_buf[1030];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1029] = exp_valid ? exp_out[1029] : encrypted_data_buf[1029];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1028] = exp_valid ? exp_out[1028] : encrypted_data_buf[1028];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1027] = exp_valid ? exp_out[1027] : encrypted_data_buf[1027];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1026] = exp_valid ? exp_out[1026] : encrypted_data_buf[1026];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1025] = exp_valid ? exp_out[1025] : encrypted_data_buf[1025];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1024] = exp_valid ? exp_out[1024] : encrypted_data_buf[1024];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1023] = exp_valid ? exp_out[1023] : encrypted_data_buf[1023];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1022] = exp_valid ? exp_out[1022] : encrypted_data_buf[1022];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1021] = exp_valid ? exp_out[1021] : encrypted_data_buf[1021];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1020] = exp_valid ? exp_out[1020] : encrypted_data_buf[1020];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1019] = exp_valid ? exp_out[1019] : encrypted_data_buf[1019];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1018] = exp_valid ? exp_out[1018] : encrypted_data_buf[1018];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1017] = exp_valid ? exp_out[1017] : encrypted_data_buf[1017];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1016] = exp_valid ? exp_out[1016] : encrypted_data_buf[1016];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1015] = exp_valid ? exp_out[1015] : encrypted_data_buf[1015];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1014] = exp_valid ? exp_out[1014] : encrypted_data_buf[1014];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1013] = exp_valid ? exp_out[1013] : encrypted_data_buf[1013];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1012] = exp_valid ? exp_out[1012] : encrypted_data_buf[1012];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1011] = exp_valid ? exp_out[1011] : encrypted_data_buf[1011];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1010] = exp_valid ? exp_out[1010] : encrypted_data_buf[1010];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1009] = exp_valid ? exp_out[1009] : encrypted_data_buf[1009];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1008] = exp_valid ? exp_out[1008] : encrypted_data_buf[1008];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1007] = exp_valid ? exp_out[1007] : encrypted_data_buf[1007];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1006] = exp_valid ? exp_out[1006] : encrypted_data_buf[1006];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1005] = exp_valid ? exp_out[1005] : encrypted_data_buf[1005];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1004] = exp_valid ? exp_out[1004] : encrypted_data_buf[1004];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1003] = exp_valid ? exp_out[1003] : encrypted_data_buf[1003];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1002] = exp_valid ? exp_out[1002] : encrypted_data_buf[1002];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1001] = exp_valid ? exp_out[1001] : encrypted_data_buf[1001];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1000] = exp_valid ? exp_out[1000] : encrypted_data_buf[1000];   // modexp_top.v(222)
    assign encrypted_data_buf_next[999] = exp_valid ? exp_out[999] : encrypted_data_buf[999];   // modexp_top.v(222)
    assign encrypted_data_buf_next[998] = exp_valid ? exp_out[998] : encrypted_data_buf[998];   // modexp_top.v(222)
    assign encrypted_data_buf_next[997] = exp_valid ? exp_out[997] : encrypted_data_buf[997];   // modexp_top.v(222)
    assign encrypted_data_buf_next[996] = exp_valid ? exp_out[996] : encrypted_data_buf[996];   // modexp_top.v(222)
    assign encrypted_data_buf_next[995] = exp_valid ? exp_out[995] : encrypted_data_buf[995];   // modexp_top.v(222)
    assign encrypted_data_buf_next[994] = exp_valid ? exp_out[994] : encrypted_data_buf[994];   // modexp_top.v(222)
    assign encrypted_data_buf_next[993] = exp_valid ? exp_out[993] : encrypted_data_buf[993];   // modexp_top.v(222)
    assign encrypted_data_buf_next[992] = exp_valid ? exp_out[992] : encrypted_data_buf[992];   // modexp_top.v(222)
    assign encrypted_data_buf_next[991] = exp_valid ? exp_out[991] : encrypted_data_buf[991];   // modexp_top.v(222)
    assign encrypted_data_buf_next[990] = exp_valid ? exp_out[990] : encrypted_data_buf[990];   // modexp_top.v(222)
    assign encrypted_data_buf_next[989] = exp_valid ? exp_out[989] : encrypted_data_buf[989];   // modexp_top.v(222)
    assign encrypted_data_buf_next[988] = exp_valid ? exp_out[988] : encrypted_data_buf[988];   // modexp_top.v(222)
    assign encrypted_data_buf_next[987] = exp_valid ? exp_out[987] : encrypted_data_buf[987];   // modexp_top.v(222)
    assign encrypted_data_buf_next[986] = exp_valid ? exp_out[986] : encrypted_data_buf[986];   // modexp_top.v(222)
    assign encrypted_data_buf_next[985] = exp_valid ? exp_out[985] : encrypted_data_buf[985];   // modexp_top.v(222)
    assign encrypted_data_buf_next[984] = exp_valid ? exp_out[984] : encrypted_data_buf[984];   // modexp_top.v(222)
    assign encrypted_data_buf_next[983] = exp_valid ? exp_out[983] : encrypted_data_buf[983];   // modexp_top.v(222)
    assign encrypted_data_buf_next[982] = exp_valid ? exp_out[982] : encrypted_data_buf[982];   // modexp_top.v(222)
    assign encrypted_data_buf_next[981] = exp_valid ? exp_out[981] : encrypted_data_buf[981];   // modexp_top.v(222)
    assign encrypted_data_buf_next[980] = exp_valid ? exp_out[980] : encrypted_data_buf[980];   // modexp_top.v(222)
    assign encrypted_data_buf_next[979] = exp_valid ? exp_out[979] : encrypted_data_buf[979];   // modexp_top.v(222)
    assign encrypted_data_buf_next[978] = exp_valid ? exp_out[978] : encrypted_data_buf[978];   // modexp_top.v(222)
    assign encrypted_data_buf_next[977] = exp_valid ? exp_out[977] : encrypted_data_buf[977];   // modexp_top.v(222)
    assign encrypted_data_buf_next[976] = exp_valid ? exp_out[976] : encrypted_data_buf[976];   // modexp_top.v(222)
    assign encrypted_data_buf_next[975] = exp_valid ? exp_out[975] : encrypted_data_buf[975];   // modexp_top.v(222)
    assign encrypted_data_buf_next[974] = exp_valid ? exp_out[974] : encrypted_data_buf[974];   // modexp_top.v(222)
    assign encrypted_data_buf_next[973] = exp_valid ? exp_out[973] : encrypted_data_buf[973];   // modexp_top.v(222)
    assign encrypted_data_buf_next[972] = exp_valid ? exp_out[972] : encrypted_data_buf[972];   // modexp_top.v(222)
    assign encrypted_data_buf_next[971] = exp_valid ? exp_out[971] : encrypted_data_buf[971];   // modexp_top.v(222)
    assign encrypted_data_buf_next[970] = exp_valid ? exp_out[970] : encrypted_data_buf[970];   // modexp_top.v(222)
    assign encrypted_data_buf_next[969] = exp_valid ? exp_out[969] : encrypted_data_buf[969];   // modexp_top.v(222)
    assign encrypted_data_buf_next[968] = exp_valid ? exp_out[968] : encrypted_data_buf[968];   // modexp_top.v(222)
    assign encrypted_data_buf_next[967] = exp_valid ? exp_out[967] : encrypted_data_buf[967];   // modexp_top.v(222)
    assign encrypted_data_buf_next[966] = exp_valid ? exp_out[966] : encrypted_data_buf[966];   // modexp_top.v(222)
    assign encrypted_data_buf_next[965] = exp_valid ? exp_out[965] : encrypted_data_buf[965];   // modexp_top.v(222)
    assign encrypted_data_buf_next[964] = exp_valid ? exp_out[964] : encrypted_data_buf[964];   // modexp_top.v(222)
    assign encrypted_data_buf_next[963] = exp_valid ? exp_out[963] : encrypted_data_buf[963];   // modexp_top.v(222)
    assign encrypted_data_buf_next[962] = exp_valid ? exp_out[962] : encrypted_data_buf[962];   // modexp_top.v(222)
    assign encrypted_data_buf_next[961] = exp_valid ? exp_out[961] : encrypted_data_buf[961];   // modexp_top.v(222)
    assign encrypted_data_buf_next[960] = exp_valid ? exp_out[960] : encrypted_data_buf[960];   // modexp_top.v(222)
    assign encrypted_data_buf_next[959] = exp_valid ? exp_out[959] : encrypted_data_buf[959];   // modexp_top.v(222)
    assign encrypted_data_buf_next[958] = exp_valid ? exp_out[958] : encrypted_data_buf[958];   // modexp_top.v(222)
    assign encrypted_data_buf_next[957] = exp_valid ? exp_out[957] : encrypted_data_buf[957];   // modexp_top.v(222)
    assign encrypted_data_buf_next[956] = exp_valid ? exp_out[956] : encrypted_data_buf[956];   // modexp_top.v(222)
    assign encrypted_data_buf_next[955] = exp_valid ? exp_out[955] : encrypted_data_buf[955];   // modexp_top.v(222)
    assign encrypted_data_buf_next[954] = exp_valid ? exp_out[954] : encrypted_data_buf[954];   // modexp_top.v(222)
    assign encrypted_data_buf_next[953] = exp_valid ? exp_out[953] : encrypted_data_buf[953];   // modexp_top.v(222)
    assign encrypted_data_buf_next[952] = exp_valid ? exp_out[952] : encrypted_data_buf[952];   // modexp_top.v(222)
    assign encrypted_data_buf_next[951] = exp_valid ? exp_out[951] : encrypted_data_buf[951];   // modexp_top.v(222)
    assign encrypted_data_buf_next[950] = exp_valid ? exp_out[950] : encrypted_data_buf[950];   // modexp_top.v(222)
    assign encrypted_data_buf_next[949] = exp_valid ? exp_out[949] : encrypted_data_buf[949];   // modexp_top.v(222)
    assign encrypted_data_buf_next[948] = exp_valid ? exp_out[948] : encrypted_data_buf[948];   // modexp_top.v(222)
    assign encrypted_data_buf_next[947] = exp_valid ? exp_out[947] : encrypted_data_buf[947];   // modexp_top.v(222)
    assign encrypted_data_buf_next[946] = exp_valid ? exp_out[946] : encrypted_data_buf[946];   // modexp_top.v(222)
    assign encrypted_data_buf_next[945] = exp_valid ? exp_out[945] : encrypted_data_buf[945];   // modexp_top.v(222)
    assign encrypted_data_buf_next[944] = exp_valid ? exp_out[944] : encrypted_data_buf[944];   // modexp_top.v(222)
    assign encrypted_data_buf_next[943] = exp_valid ? exp_out[943] : encrypted_data_buf[943];   // modexp_top.v(222)
    assign encrypted_data_buf_next[942] = exp_valid ? exp_out[942] : encrypted_data_buf[942];   // modexp_top.v(222)
    assign encrypted_data_buf_next[941] = exp_valid ? exp_out[941] : encrypted_data_buf[941];   // modexp_top.v(222)
    assign encrypted_data_buf_next[940] = exp_valid ? exp_out[940] : encrypted_data_buf[940];   // modexp_top.v(222)
    assign encrypted_data_buf_next[939] = exp_valid ? exp_out[939] : encrypted_data_buf[939];   // modexp_top.v(222)
    assign encrypted_data_buf_next[938] = exp_valid ? exp_out[938] : encrypted_data_buf[938];   // modexp_top.v(222)
    assign encrypted_data_buf_next[937] = exp_valid ? exp_out[937] : encrypted_data_buf[937];   // modexp_top.v(222)
    assign encrypted_data_buf_next[936] = exp_valid ? exp_out[936] : encrypted_data_buf[936];   // modexp_top.v(222)
    assign encrypted_data_buf_next[935] = exp_valid ? exp_out[935] : encrypted_data_buf[935];   // modexp_top.v(222)
    assign encrypted_data_buf_next[934] = exp_valid ? exp_out[934] : encrypted_data_buf[934];   // modexp_top.v(222)
    assign encrypted_data_buf_next[933] = exp_valid ? exp_out[933] : encrypted_data_buf[933];   // modexp_top.v(222)
    assign encrypted_data_buf_next[932] = exp_valid ? exp_out[932] : encrypted_data_buf[932];   // modexp_top.v(222)
    assign encrypted_data_buf_next[931] = exp_valid ? exp_out[931] : encrypted_data_buf[931];   // modexp_top.v(222)
    assign encrypted_data_buf_next[930] = exp_valid ? exp_out[930] : encrypted_data_buf[930];   // modexp_top.v(222)
    assign encrypted_data_buf_next[929] = exp_valid ? exp_out[929] : encrypted_data_buf[929];   // modexp_top.v(222)
    assign encrypted_data_buf_next[928] = exp_valid ? exp_out[928] : encrypted_data_buf[928];   // modexp_top.v(222)
    assign encrypted_data_buf_next[927] = exp_valid ? exp_out[927] : encrypted_data_buf[927];   // modexp_top.v(222)
    assign encrypted_data_buf_next[926] = exp_valid ? exp_out[926] : encrypted_data_buf[926];   // modexp_top.v(222)
    assign encrypted_data_buf_next[925] = exp_valid ? exp_out[925] : encrypted_data_buf[925];   // modexp_top.v(222)
    assign encrypted_data_buf_next[924] = exp_valid ? exp_out[924] : encrypted_data_buf[924];   // modexp_top.v(222)
    assign encrypted_data_buf_next[923] = exp_valid ? exp_out[923] : encrypted_data_buf[923];   // modexp_top.v(222)
    assign encrypted_data_buf_next[922] = exp_valid ? exp_out[922] : encrypted_data_buf[922];   // modexp_top.v(222)
    assign encrypted_data_buf_next[921] = exp_valid ? exp_out[921] : encrypted_data_buf[921];   // modexp_top.v(222)
    assign encrypted_data_buf_next[920] = exp_valid ? exp_out[920] : encrypted_data_buf[920];   // modexp_top.v(222)
    assign encrypted_data_buf_next[919] = exp_valid ? exp_out[919] : encrypted_data_buf[919];   // modexp_top.v(222)
    assign encrypted_data_buf_next[918] = exp_valid ? exp_out[918] : encrypted_data_buf[918];   // modexp_top.v(222)
    assign encrypted_data_buf_next[917] = exp_valid ? exp_out[917] : encrypted_data_buf[917];   // modexp_top.v(222)
    assign encrypted_data_buf_next[916] = exp_valid ? exp_out[916] : encrypted_data_buf[916];   // modexp_top.v(222)
    assign encrypted_data_buf_next[915] = exp_valid ? exp_out[915] : encrypted_data_buf[915];   // modexp_top.v(222)
    assign encrypted_data_buf_next[914] = exp_valid ? exp_out[914] : encrypted_data_buf[914];   // modexp_top.v(222)
    assign encrypted_data_buf_next[913] = exp_valid ? exp_out[913] : encrypted_data_buf[913];   // modexp_top.v(222)
    assign encrypted_data_buf_next[912] = exp_valid ? exp_out[912] : encrypted_data_buf[912];   // modexp_top.v(222)
    assign encrypted_data_buf_next[911] = exp_valid ? exp_out[911] : encrypted_data_buf[911];   // modexp_top.v(222)
    assign encrypted_data_buf_next[910] = exp_valid ? exp_out[910] : encrypted_data_buf[910];   // modexp_top.v(222)
    assign encrypted_data_buf_next[909] = exp_valid ? exp_out[909] : encrypted_data_buf[909];   // modexp_top.v(222)
    assign encrypted_data_buf_next[908] = exp_valid ? exp_out[908] : encrypted_data_buf[908];   // modexp_top.v(222)
    assign encrypted_data_buf_next[907] = exp_valid ? exp_out[907] : encrypted_data_buf[907];   // modexp_top.v(222)
    assign encrypted_data_buf_next[906] = exp_valid ? exp_out[906] : encrypted_data_buf[906];   // modexp_top.v(222)
    assign encrypted_data_buf_next[905] = exp_valid ? exp_out[905] : encrypted_data_buf[905];   // modexp_top.v(222)
    assign encrypted_data_buf_next[904] = exp_valid ? exp_out[904] : encrypted_data_buf[904];   // modexp_top.v(222)
    assign encrypted_data_buf_next[903] = exp_valid ? exp_out[903] : encrypted_data_buf[903];   // modexp_top.v(222)
    assign encrypted_data_buf_next[902] = exp_valid ? exp_out[902] : encrypted_data_buf[902];   // modexp_top.v(222)
    assign encrypted_data_buf_next[901] = exp_valid ? exp_out[901] : encrypted_data_buf[901];   // modexp_top.v(222)
    assign encrypted_data_buf_next[900] = exp_valid ? exp_out[900] : encrypted_data_buf[900];   // modexp_top.v(222)
    assign encrypted_data_buf_next[899] = exp_valid ? exp_out[899] : encrypted_data_buf[899];   // modexp_top.v(222)
    assign encrypted_data_buf_next[898] = exp_valid ? exp_out[898] : encrypted_data_buf[898];   // modexp_top.v(222)
    assign encrypted_data_buf_next[897] = exp_valid ? exp_out[897] : encrypted_data_buf[897];   // modexp_top.v(222)
    assign encrypted_data_buf_next[896] = exp_valid ? exp_out[896] : encrypted_data_buf[896];   // modexp_top.v(222)
    assign encrypted_data_buf_next[895] = exp_valid ? exp_out[895] : encrypted_data_buf[895];   // modexp_top.v(222)
    assign encrypted_data_buf_next[894] = exp_valid ? exp_out[894] : encrypted_data_buf[894];   // modexp_top.v(222)
    assign encrypted_data_buf_next[893] = exp_valid ? exp_out[893] : encrypted_data_buf[893];   // modexp_top.v(222)
    assign encrypted_data_buf_next[892] = exp_valid ? exp_out[892] : encrypted_data_buf[892];   // modexp_top.v(222)
    assign encrypted_data_buf_next[891] = exp_valid ? exp_out[891] : encrypted_data_buf[891];   // modexp_top.v(222)
    assign encrypted_data_buf_next[890] = exp_valid ? exp_out[890] : encrypted_data_buf[890];   // modexp_top.v(222)
    assign encrypted_data_buf_next[889] = exp_valid ? exp_out[889] : encrypted_data_buf[889];   // modexp_top.v(222)
    assign encrypted_data_buf_next[888] = exp_valid ? exp_out[888] : encrypted_data_buf[888];   // modexp_top.v(222)
    assign encrypted_data_buf_next[887] = exp_valid ? exp_out[887] : encrypted_data_buf[887];   // modexp_top.v(222)
    assign encrypted_data_buf_next[886] = exp_valid ? exp_out[886] : encrypted_data_buf[886];   // modexp_top.v(222)
    assign encrypted_data_buf_next[885] = exp_valid ? exp_out[885] : encrypted_data_buf[885];   // modexp_top.v(222)
    assign encrypted_data_buf_next[884] = exp_valid ? exp_out[884] : encrypted_data_buf[884];   // modexp_top.v(222)
    assign encrypted_data_buf_next[883] = exp_valid ? exp_out[883] : encrypted_data_buf[883];   // modexp_top.v(222)
    assign encrypted_data_buf_next[882] = exp_valid ? exp_out[882] : encrypted_data_buf[882];   // modexp_top.v(222)
    assign encrypted_data_buf_next[881] = exp_valid ? exp_out[881] : encrypted_data_buf[881];   // modexp_top.v(222)
    assign encrypted_data_buf_next[880] = exp_valid ? exp_out[880] : encrypted_data_buf[880];   // modexp_top.v(222)
    assign encrypted_data_buf_next[879] = exp_valid ? exp_out[879] : encrypted_data_buf[879];   // modexp_top.v(222)
    assign encrypted_data_buf_next[878] = exp_valid ? exp_out[878] : encrypted_data_buf[878];   // modexp_top.v(222)
    assign encrypted_data_buf_next[877] = exp_valid ? exp_out[877] : encrypted_data_buf[877];   // modexp_top.v(222)
    assign encrypted_data_buf_next[876] = exp_valid ? exp_out[876] : encrypted_data_buf[876];   // modexp_top.v(222)
    assign encrypted_data_buf_next[875] = exp_valid ? exp_out[875] : encrypted_data_buf[875];   // modexp_top.v(222)
    assign encrypted_data_buf_next[874] = exp_valid ? exp_out[874] : encrypted_data_buf[874];   // modexp_top.v(222)
    assign encrypted_data_buf_next[873] = exp_valid ? exp_out[873] : encrypted_data_buf[873];   // modexp_top.v(222)
    assign encrypted_data_buf_next[872] = exp_valid ? exp_out[872] : encrypted_data_buf[872];   // modexp_top.v(222)
    assign encrypted_data_buf_next[871] = exp_valid ? exp_out[871] : encrypted_data_buf[871];   // modexp_top.v(222)
    assign encrypted_data_buf_next[870] = exp_valid ? exp_out[870] : encrypted_data_buf[870];   // modexp_top.v(222)
    assign encrypted_data_buf_next[869] = exp_valid ? exp_out[869] : encrypted_data_buf[869];   // modexp_top.v(222)
    assign encrypted_data_buf_next[868] = exp_valid ? exp_out[868] : encrypted_data_buf[868];   // modexp_top.v(222)
    assign encrypted_data_buf_next[867] = exp_valid ? exp_out[867] : encrypted_data_buf[867];   // modexp_top.v(222)
    assign encrypted_data_buf_next[866] = exp_valid ? exp_out[866] : encrypted_data_buf[866];   // modexp_top.v(222)
    assign encrypted_data_buf_next[865] = exp_valid ? exp_out[865] : encrypted_data_buf[865];   // modexp_top.v(222)
    assign encrypted_data_buf_next[864] = exp_valid ? exp_out[864] : encrypted_data_buf[864];   // modexp_top.v(222)
    assign encrypted_data_buf_next[863] = exp_valid ? exp_out[863] : encrypted_data_buf[863];   // modexp_top.v(222)
    assign encrypted_data_buf_next[862] = exp_valid ? exp_out[862] : encrypted_data_buf[862];   // modexp_top.v(222)
    assign encrypted_data_buf_next[861] = exp_valid ? exp_out[861] : encrypted_data_buf[861];   // modexp_top.v(222)
    assign encrypted_data_buf_next[860] = exp_valid ? exp_out[860] : encrypted_data_buf[860];   // modexp_top.v(222)
    assign encrypted_data_buf_next[859] = exp_valid ? exp_out[859] : encrypted_data_buf[859];   // modexp_top.v(222)
    assign encrypted_data_buf_next[858] = exp_valid ? exp_out[858] : encrypted_data_buf[858];   // modexp_top.v(222)
    assign encrypted_data_buf_next[857] = exp_valid ? exp_out[857] : encrypted_data_buf[857];   // modexp_top.v(222)
    assign encrypted_data_buf_next[856] = exp_valid ? exp_out[856] : encrypted_data_buf[856];   // modexp_top.v(222)
    assign encrypted_data_buf_next[855] = exp_valid ? exp_out[855] : encrypted_data_buf[855];   // modexp_top.v(222)
    assign encrypted_data_buf_next[854] = exp_valid ? exp_out[854] : encrypted_data_buf[854];   // modexp_top.v(222)
    assign encrypted_data_buf_next[853] = exp_valid ? exp_out[853] : encrypted_data_buf[853];   // modexp_top.v(222)
    assign encrypted_data_buf_next[852] = exp_valid ? exp_out[852] : encrypted_data_buf[852];   // modexp_top.v(222)
    assign encrypted_data_buf_next[851] = exp_valid ? exp_out[851] : encrypted_data_buf[851];   // modexp_top.v(222)
    assign encrypted_data_buf_next[850] = exp_valid ? exp_out[850] : encrypted_data_buf[850];   // modexp_top.v(222)
    assign encrypted_data_buf_next[849] = exp_valid ? exp_out[849] : encrypted_data_buf[849];   // modexp_top.v(222)
    assign encrypted_data_buf_next[848] = exp_valid ? exp_out[848] : encrypted_data_buf[848];   // modexp_top.v(222)
    assign encrypted_data_buf_next[847] = exp_valid ? exp_out[847] : encrypted_data_buf[847];   // modexp_top.v(222)
    assign encrypted_data_buf_next[846] = exp_valid ? exp_out[846] : encrypted_data_buf[846];   // modexp_top.v(222)
    assign encrypted_data_buf_next[845] = exp_valid ? exp_out[845] : encrypted_data_buf[845];   // modexp_top.v(222)
    assign encrypted_data_buf_next[844] = exp_valid ? exp_out[844] : encrypted_data_buf[844];   // modexp_top.v(222)
    assign encrypted_data_buf_next[843] = exp_valid ? exp_out[843] : encrypted_data_buf[843];   // modexp_top.v(222)
    assign encrypted_data_buf_next[842] = exp_valid ? exp_out[842] : encrypted_data_buf[842];   // modexp_top.v(222)
    assign encrypted_data_buf_next[841] = exp_valid ? exp_out[841] : encrypted_data_buf[841];   // modexp_top.v(222)
    assign encrypted_data_buf_next[840] = exp_valid ? exp_out[840] : encrypted_data_buf[840];   // modexp_top.v(222)
    assign encrypted_data_buf_next[839] = exp_valid ? exp_out[839] : encrypted_data_buf[839];   // modexp_top.v(222)
    assign encrypted_data_buf_next[838] = exp_valid ? exp_out[838] : encrypted_data_buf[838];   // modexp_top.v(222)
    assign encrypted_data_buf_next[837] = exp_valid ? exp_out[837] : encrypted_data_buf[837];   // modexp_top.v(222)
    assign encrypted_data_buf_next[836] = exp_valid ? exp_out[836] : encrypted_data_buf[836];   // modexp_top.v(222)
    assign encrypted_data_buf_next[835] = exp_valid ? exp_out[835] : encrypted_data_buf[835];   // modexp_top.v(222)
    assign encrypted_data_buf_next[834] = exp_valid ? exp_out[834] : encrypted_data_buf[834];   // modexp_top.v(222)
    assign encrypted_data_buf_next[833] = exp_valid ? exp_out[833] : encrypted_data_buf[833];   // modexp_top.v(222)
    assign encrypted_data_buf_next[832] = exp_valid ? exp_out[832] : encrypted_data_buf[832];   // modexp_top.v(222)
    assign encrypted_data_buf_next[831] = exp_valid ? exp_out[831] : encrypted_data_buf[831];   // modexp_top.v(222)
    assign encrypted_data_buf_next[830] = exp_valid ? exp_out[830] : encrypted_data_buf[830];   // modexp_top.v(222)
    assign encrypted_data_buf_next[829] = exp_valid ? exp_out[829] : encrypted_data_buf[829];   // modexp_top.v(222)
    assign encrypted_data_buf_next[828] = exp_valid ? exp_out[828] : encrypted_data_buf[828];   // modexp_top.v(222)
    assign encrypted_data_buf_next[827] = exp_valid ? exp_out[827] : encrypted_data_buf[827];   // modexp_top.v(222)
    assign encrypted_data_buf_next[826] = exp_valid ? exp_out[826] : encrypted_data_buf[826];   // modexp_top.v(222)
    assign encrypted_data_buf_next[825] = exp_valid ? exp_out[825] : encrypted_data_buf[825];   // modexp_top.v(222)
    assign encrypted_data_buf_next[824] = exp_valid ? exp_out[824] : encrypted_data_buf[824];   // modexp_top.v(222)
    assign encrypted_data_buf_next[823] = exp_valid ? exp_out[823] : encrypted_data_buf[823];   // modexp_top.v(222)
    assign encrypted_data_buf_next[822] = exp_valid ? exp_out[822] : encrypted_data_buf[822];   // modexp_top.v(222)
    assign encrypted_data_buf_next[821] = exp_valid ? exp_out[821] : encrypted_data_buf[821];   // modexp_top.v(222)
    assign encrypted_data_buf_next[820] = exp_valid ? exp_out[820] : encrypted_data_buf[820];   // modexp_top.v(222)
    assign encrypted_data_buf_next[819] = exp_valid ? exp_out[819] : encrypted_data_buf[819];   // modexp_top.v(222)
    assign encrypted_data_buf_next[818] = exp_valid ? exp_out[818] : encrypted_data_buf[818];   // modexp_top.v(222)
    assign encrypted_data_buf_next[817] = exp_valid ? exp_out[817] : encrypted_data_buf[817];   // modexp_top.v(222)
    assign encrypted_data_buf_next[816] = exp_valid ? exp_out[816] : encrypted_data_buf[816];   // modexp_top.v(222)
    assign encrypted_data_buf_next[815] = exp_valid ? exp_out[815] : encrypted_data_buf[815];   // modexp_top.v(222)
    assign encrypted_data_buf_next[814] = exp_valid ? exp_out[814] : encrypted_data_buf[814];   // modexp_top.v(222)
    assign encrypted_data_buf_next[813] = exp_valid ? exp_out[813] : encrypted_data_buf[813];   // modexp_top.v(222)
    assign encrypted_data_buf_next[812] = exp_valid ? exp_out[812] : encrypted_data_buf[812];   // modexp_top.v(222)
    assign encrypted_data_buf_next[811] = exp_valid ? exp_out[811] : encrypted_data_buf[811];   // modexp_top.v(222)
    assign encrypted_data_buf_next[810] = exp_valid ? exp_out[810] : encrypted_data_buf[810];   // modexp_top.v(222)
    assign encrypted_data_buf_next[809] = exp_valid ? exp_out[809] : encrypted_data_buf[809];   // modexp_top.v(222)
    assign encrypted_data_buf_next[808] = exp_valid ? exp_out[808] : encrypted_data_buf[808];   // modexp_top.v(222)
    assign encrypted_data_buf_next[807] = exp_valid ? exp_out[807] : encrypted_data_buf[807];   // modexp_top.v(222)
    assign encrypted_data_buf_next[806] = exp_valid ? exp_out[806] : encrypted_data_buf[806];   // modexp_top.v(222)
    assign encrypted_data_buf_next[805] = exp_valid ? exp_out[805] : encrypted_data_buf[805];   // modexp_top.v(222)
    assign encrypted_data_buf_next[804] = exp_valid ? exp_out[804] : encrypted_data_buf[804];   // modexp_top.v(222)
    assign encrypted_data_buf_next[803] = exp_valid ? exp_out[803] : encrypted_data_buf[803];   // modexp_top.v(222)
    assign encrypted_data_buf_next[802] = exp_valid ? exp_out[802] : encrypted_data_buf[802];   // modexp_top.v(222)
    assign encrypted_data_buf_next[801] = exp_valid ? exp_out[801] : encrypted_data_buf[801];   // modexp_top.v(222)
    assign encrypted_data_buf_next[800] = exp_valid ? exp_out[800] : encrypted_data_buf[800];   // modexp_top.v(222)
    assign encrypted_data_buf_next[799] = exp_valid ? exp_out[799] : encrypted_data_buf[799];   // modexp_top.v(222)
    assign encrypted_data_buf_next[798] = exp_valid ? exp_out[798] : encrypted_data_buf[798];   // modexp_top.v(222)
    assign encrypted_data_buf_next[797] = exp_valid ? exp_out[797] : encrypted_data_buf[797];   // modexp_top.v(222)
    assign encrypted_data_buf_next[796] = exp_valid ? exp_out[796] : encrypted_data_buf[796];   // modexp_top.v(222)
    assign encrypted_data_buf_next[795] = exp_valid ? exp_out[795] : encrypted_data_buf[795];   // modexp_top.v(222)
    assign encrypted_data_buf_next[794] = exp_valid ? exp_out[794] : encrypted_data_buf[794];   // modexp_top.v(222)
    assign encrypted_data_buf_next[793] = exp_valid ? exp_out[793] : encrypted_data_buf[793];   // modexp_top.v(222)
    assign encrypted_data_buf_next[792] = exp_valid ? exp_out[792] : encrypted_data_buf[792];   // modexp_top.v(222)
    assign encrypted_data_buf_next[791] = exp_valid ? exp_out[791] : encrypted_data_buf[791];   // modexp_top.v(222)
    assign encrypted_data_buf_next[790] = exp_valid ? exp_out[790] : encrypted_data_buf[790];   // modexp_top.v(222)
    assign encrypted_data_buf_next[789] = exp_valid ? exp_out[789] : encrypted_data_buf[789];   // modexp_top.v(222)
    assign encrypted_data_buf_next[788] = exp_valid ? exp_out[788] : encrypted_data_buf[788];   // modexp_top.v(222)
    assign encrypted_data_buf_next[787] = exp_valid ? exp_out[787] : encrypted_data_buf[787];   // modexp_top.v(222)
    assign encrypted_data_buf_next[786] = exp_valid ? exp_out[786] : encrypted_data_buf[786];   // modexp_top.v(222)
    assign encrypted_data_buf_next[785] = exp_valid ? exp_out[785] : encrypted_data_buf[785];   // modexp_top.v(222)
    assign encrypted_data_buf_next[784] = exp_valid ? exp_out[784] : encrypted_data_buf[784];   // modexp_top.v(222)
    assign encrypted_data_buf_next[783] = exp_valid ? exp_out[783] : encrypted_data_buf[783];   // modexp_top.v(222)
    assign encrypted_data_buf_next[782] = exp_valid ? exp_out[782] : encrypted_data_buf[782];   // modexp_top.v(222)
    assign encrypted_data_buf_next[781] = exp_valid ? exp_out[781] : encrypted_data_buf[781];   // modexp_top.v(222)
    assign encrypted_data_buf_next[780] = exp_valid ? exp_out[780] : encrypted_data_buf[780];   // modexp_top.v(222)
    assign encrypted_data_buf_next[779] = exp_valid ? exp_out[779] : encrypted_data_buf[779];   // modexp_top.v(222)
    assign encrypted_data_buf_next[778] = exp_valid ? exp_out[778] : encrypted_data_buf[778];   // modexp_top.v(222)
    assign encrypted_data_buf_next[777] = exp_valid ? exp_out[777] : encrypted_data_buf[777];   // modexp_top.v(222)
    assign encrypted_data_buf_next[776] = exp_valid ? exp_out[776] : encrypted_data_buf[776];   // modexp_top.v(222)
    assign encrypted_data_buf_next[775] = exp_valid ? exp_out[775] : encrypted_data_buf[775];   // modexp_top.v(222)
    assign encrypted_data_buf_next[774] = exp_valid ? exp_out[774] : encrypted_data_buf[774];   // modexp_top.v(222)
    assign encrypted_data_buf_next[773] = exp_valid ? exp_out[773] : encrypted_data_buf[773];   // modexp_top.v(222)
    assign encrypted_data_buf_next[772] = exp_valid ? exp_out[772] : encrypted_data_buf[772];   // modexp_top.v(222)
    assign encrypted_data_buf_next[771] = exp_valid ? exp_out[771] : encrypted_data_buf[771];   // modexp_top.v(222)
    assign encrypted_data_buf_next[770] = exp_valid ? exp_out[770] : encrypted_data_buf[770];   // modexp_top.v(222)
    assign encrypted_data_buf_next[769] = exp_valid ? exp_out[769] : encrypted_data_buf[769];   // modexp_top.v(222)
    assign encrypted_data_buf_next[768] = exp_valid ? exp_out[768] : encrypted_data_buf[768];   // modexp_top.v(222)
    assign encrypted_data_buf_next[767] = exp_valid ? exp_out[767] : encrypted_data_buf[767];   // modexp_top.v(222)
    assign encrypted_data_buf_next[766] = exp_valid ? exp_out[766] : encrypted_data_buf[766];   // modexp_top.v(222)
    assign encrypted_data_buf_next[765] = exp_valid ? exp_out[765] : encrypted_data_buf[765];   // modexp_top.v(222)
    assign encrypted_data_buf_next[764] = exp_valid ? exp_out[764] : encrypted_data_buf[764];   // modexp_top.v(222)
    assign encrypted_data_buf_next[763] = exp_valid ? exp_out[763] : encrypted_data_buf[763];   // modexp_top.v(222)
    assign encrypted_data_buf_next[762] = exp_valid ? exp_out[762] : encrypted_data_buf[762];   // modexp_top.v(222)
    assign encrypted_data_buf_next[761] = exp_valid ? exp_out[761] : encrypted_data_buf[761];   // modexp_top.v(222)
    assign encrypted_data_buf_next[760] = exp_valid ? exp_out[760] : encrypted_data_buf[760];   // modexp_top.v(222)
    assign encrypted_data_buf_next[759] = exp_valid ? exp_out[759] : encrypted_data_buf[759];   // modexp_top.v(222)
    assign encrypted_data_buf_next[758] = exp_valid ? exp_out[758] : encrypted_data_buf[758];   // modexp_top.v(222)
    assign encrypted_data_buf_next[757] = exp_valid ? exp_out[757] : encrypted_data_buf[757];   // modexp_top.v(222)
    assign encrypted_data_buf_next[756] = exp_valid ? exp_out[756] : encrypted_data_buf[756];   // modexp_top.v(222)
    assign encrypted_data_buf_next[755] = exp_valid ? exp_out[755] : encrypted_data_buf[755];   // modexp_top.v(222)
    assign encrypted_data_buf_next[754] = exp_valid ? exp_out[754] : encrypted_data_buf[754];   // modexp_top.v(222)
    assign encrypted_data_buf_next[753] = exp_valid ? exp_out[753] : encrypted_data_buf[753];   // modexp_top.v(222)
    assign encrypted_data_buf_next[752] = exp_valid ? exp_out[752] : encrypted_data_buf[752];   // modexp_top.v(222)
    assign encrypted_data_buf_next[751] = exp_valid ? exp_out[751] : encrypted_data_buf[751];   // modexp_top.v(222)
    assign encrypted_data_buf_next[750] = exp_valid ? exp_out[750] : encrypted_data_buf[750];   // modexp_top.v(222)
    assign encrypted_data_buf_next[749] = exp_valid ? exp_out[749] : encrypted_data_buf[749];   // modexp_top.v(222)
    assign encrypted_data_buf_next[748] = exp_valid ? exp_out[748] : encrypted_data_buf[748];   // modexp_top.v(222)
    assign encrypted_data_buf_next[747] = exp_valid ? exp_out[747] : encrypted_data_buf[747];   // modexp_top.v(222)
    assign encrypted_data_buf_next[746] = exp_valid ? exp_out[746] : encrypted_data_buf[746];   // modexp_top.v(222)
    assign encrypted_data_buf_next[745] = exp_valid ? exp_out[745] : encrypted_data_buf[745];   // modexp_top.v(222)
    assign encrypted_data_buf_next[744] = exp_valid ? exp_out[744] : encrypted_data_buf[744];   // modexp_top.v(222)
    assign encrypted_data_buf_next[743] = exp_valid ? exp_out[743] : encrypted_data_buf[743];   // modexp_top.v(222)
    assign encrypted_data_buf_next[742] = exp_valid ? exp_out[742] : encrypted_data_buf[742];   // modexp_top.v(222)
    assign encrypted_data_buf_next[741] = exp_valid ? exp_out[741] : encrypted_data_buf[741];   // modexp_top.v(222)
    assign encrypted_data_buf_next[740] = exp_valid ? exp_out[740] : encrypted_data_buf[740];   // modexp_top.v(222)
    assign encrypted_data_buf_next[739] = exp_valid ? exp_out[739] : encrypted_data_buf[739];   // modexp_top.v(222)
    assign encrypted_data_buf_next[738] = exp_valid ? exp_out[738] : encrypted_data_buf[738];   // modexp_top.v(222)
    assign encrypted_data_buf_next[737] = exp_valid ? exp_out[737] : encrypted_data_buf[737];   // modexp_top.v(222)
    assign encrypted_data_buf_next[736] = exp_valid ? exp_out[736] : encrypted_data_buf[736];   // modexp_top.v(222)
    assign encrypted_data_buf_next[735] = exp_valid ? exp_out[735] : encrypted_data_buf[735];   // modexp_top.v(222)
    assign encrypted_data_buf_next[734] = exp_valid ? exp_out[734] : encrypted_data_buf[734];   // modexp_top.v(222)
    assign encrypted_data_buf_next[733] = exp_valid ? exp_out[733] : encrypted_data_buf[733];   // modexp_top.v(222)
    assign encrypted_data_buf_next[732] = exp_valid ? exp_out[732] : encrypted_data_buf[732];   // modexp_top.v(222)
    assign encrypted_data_buf_next[731] = exp_valid ? exp_out[731] : encrypted_data_buf[731];   // modexp_top.v(222)
    assign encrypted_data_buf_next[730] = exp_valid ? exp_out[730] : encrypted_data_buf[730];   // modexp_top.v(222)
    assign encrypted_data_buf_next[729] = exp_valid ? exp_out[729] : encrypted_data_buf[729];   // modexp_top.v(222)
    assign encrypted_data_buf_next[728] = exp_valid ? exp_out[728] : encrypted_data_buf[728];   // modexp_top.v(222)
    assign encrypted_data_buf_next[727] = exp_valid ? exp_out[727] : encrypted_data_buf[727];   // modexp_top.v(222)
    assign encrypted_data_buf_next[726] = exp_valid ? exp_out[726] : encrypted_data_buf[726];   // modexp_top.v(222)
    assign encrypted_data_buf_next[725] = exp_valid ? exp_out[725] : encrypted_data_buf[725];   // modexp_top.v(222)
    assign encrypted_data_buf_next[724] = exp_valid ? exp_out[724] : encrypted_data_buf[724];   // modexp_top.v(222)
    assign encrypted_data_buf_next[723] = exp_valid ? exp_out[723] : encrypted_data_buf[723];   // modexp_top.v(222)
    assign encrypted_data_buf_next[722] = exp_valid ? exp_out[722] : encrypted_data_buf[722];   // modexp_top.v(222)
    assign encrypted_data_buf_next[721] = exp_valid ? exp_out[721] : encrypted_data_buf[721];   // modexp_top.v(222)
    assign encrypted_data_buf_next[720] = exp_valid ? exp_out[720] : encrypted_data_buf[720];   // modexp_top.v(222)
    assign encrypted_data_buf_next[719] = exp_valid ? exp_out[719] : encrypted_data_buf[719];   // modexp_top.v(222)
    assign encrypted_data_buf_next[718] = exp_valid ? exp_out[718] : encrypted_data_buf[718];   // modexp_top.v(222)
    assign encrypted_data_buf_next[717] = exp_valid ? exp_out[717] : encrypted_data_buf[717];   // modexp_top.v(222)
    assign encrypted_data_buf_next[716] = exp_valid ? exp_out[716] : encrypted_data_buf[716];   // modexp_top.v(222)
    assign encrypted_data_buf_next[715] = exp_valid ? exp_out[715] : encrypted_data_buf[715];   // modexp_top.v(222)
    assign encrypted_data_buf_next[714] = exp_valid ? exp_out[714] : encrypted_data_buf[714];   // modexp_top.v(222)
    assign encrypted_data_buf_next[713] = exp_valid ? exp_out[713] : encrypted_data_buf[713];   // modexp_top.v(222)
    assign encrypted_data_buf_next[712] = exp_valid ? exp_out[712] : encrypted_data_buf[712];   // modexp_top.v(222)
    assign encrypted_data_buf_next[711] = exp_valid ? exp_out[711] : encrypted_data_buf[711];   // modexp_top.v(222)
    assign encrypted_data_buf_next[710] = exp_valid ? exp_out[710] : encrypted_data_buf[710];   // modexp_top.v(222)
    assign encrypted_data_buf_next[709] = exp_valid ? exp_out[709] : encrypted_data_buf[709];   // modexp_top.v(222)
    assign encrypted_data_buf_next[708] = exp_valid ? exp_out[708] : encrypted_data_buf[708];   // modexp_top.v(222)
    assign encrypted_data_buf_next[707] = exp_valid ? exp_out[707] : encrypted_data_buf[707];   // modexp_top.v(222)
    assign encrypted_data_buf_next[706] = exp_valid ? exp_out[706] : encrypted_data_buf[706];   // modexp_top.v(222)
    assign encrypted_data_buf_next[705] = exp_valid ? exp_out[705] : encrypted_data_buf[705];   // modexp_top.v(222)
    assign encrypted_data_buf_next[704] = exp_valid ? exp_out[704] : encrypted_data_buf[704];   // modexp_top.v(222)
    assign encrypted_data_buf_next[703] = exp_valid ? exp_out[703] : encrypted_data_buf[703];   // modexp_top.v(222)
    assign encrypted_data_buf_next[702] = exp_valid ? exp_out[702] : encrypted_data_buf[702];   // modexp_top.v(222)
    assign encrypted_data_buf_next[701] = exp_valid ? exp_out[701] : encrypted_data_buf[701];   // modexp_top.v(222)
    assign encrypted_data_buf_next[700] = exp_valid ? exp_out[700] : encrypted_data_buf[700];   // modexp_top.v(222)
    assign encrypted_data_buf_next[699] = exp_valid ? exp_out[699] : encrypted_data_buf[699];   // modexp_top.v(222)
    assign encrypted_data_buf_next[698] = exp_valid ? exp_out[698] : encrypted_data_buf[698];   // modexp_top.v(222)
    assign encrypted_data_buf_next[697] = exp_valid ? exp_out[697] : encrypted_data_buf[697];   // modexp_top.v(222)
    assign encrypted_data_buf_next[696] = exp_valid ? exp_out[696] : encrypted_data_buf[696];   // modexp_top.v(222)
    assign encrypted_data_buf_next[695] = exp_valid ? exp_out[695] : encrypted_data_buf[695];   // modexp_top.v(222)
    assign encrypted_data_buf_next[694] = exp_valid ? exp_out[694] : encrypted_data_buf[694];   // modexp_top.v(222)
    assign encrypted_data_buf_next[693] = exp_valid ? exp_out[693] : encrypted_data_buf[693];   // modexp_top.v(222)
    assign encrypted_data_buf_next[692] = exp_valid ? exp_out[692] : encrypted_data_buf[692];   // modexp_top.v(222)
    assign encrypted_data_buf_next[691] = exp_valid ? exp_out[691] : encrypted_data_buf[691];   // modexp_top.v(222)
    assign encrypted_data_buf_next[690] = exp_valid ? exp_out[690] : encrypted_data_buf[690];   // modexp_top.v(222)
    assign encrypted_data_buf_next[689] = exp_valid ? exp_out[689] : encrypted_data_buf[689];   // modexp_top.v(222)
    assign encrypted_data_buf_next[688] = exp_valid ? exp_out[688] : encrypted_data_buf[688];   // modexp_top.v(222)
    assign encrypted_data_buf_next[687] = exp_valid ? exp_out[687] : encrypted_data_buf[687];   // modexp_top.v(222)
    assign encrypted_data_buf_next[686] = exp_valid ? exp_out[686] : encrypted_data_buf[686];   // modexp_top.v(222)
    assign encrypted_data_buf_next[685] = exp_valid ? exp_out[685] : encrypted_data_buf[685];   // modexp_top.v(222)
    assign encrypted_data_buf_next[684] = exp_valid ? exp_out[684] : encrypted_data_buf[684];   // modexp_top.v(222)
    assign encrypted_data_buf_next[683] = exp_valid ? exp_out[683] : encrypted_data_buf[683];   // modexp_top.v(222)
    assign encrypted_data_buf_next[682] = exp_valid ? exp_out[682] : encrypted_data_buf[682];   // modexp_top.v(222)
    assign encrypted_data_buf_next[681] = exp_valid ? exp_out[681] : encrypted_data_buf[681];   // modexp_top.v(222)
    assign encrypted_data_buf_next[680] = exp_valid ? exp_out[680] : encrypted_data_buf[680];   // modexp_top.v(222)
    assign encrypted_data_buf_next[679] = exp_valid ? exp_out[679] : encrypted_data_buf[679];   // modexp_top.v(222)
    assign encrypted_data_buf_next[678] = exp_valid ? exp_out[678] : encrypted_data_buf[678];   // modexp_top.v(222)
    assign encrypted_data_buf_next[677] = exp_valid ? exp_out[677] : encrypted_data_buf[677];   // modexp_top.v(222)
    assign encrypted_data_buf_next[676] = exp_valid ? exp_out[676] : encrypted_data_buf[676];   // modexp_top.v(222)
    assign encrypted_data_buf_next[675] = exp_valid ? exp_out[675] : encrypted_data_buf[675];   // modexp_top.v(222)
    assign encrypted_data_buf_next[674] = exp_valid ? exp_out[674] : encrypted_data_buf[674];   // modexp_top.v(222)
    assign encrypted_data_buf_next[673] = exp_valid ? exp_out[673] : encrypted_data_buf[673];   // modexp_top.v(222)
    assign encrypted_data_buf_next[672] = exp_valid ? exp_out[672] : encrypted_data_buf[672];   // modexp_top.v(222)
    assign encrypted_data_buf_next[671] = exp_valid ? exp_out[671] : encrypted_data_buf[671];   // modexp_top.v(222)
    assign encrypted_data_buf_next[670] = exp_valid ? exp_out[670] : encrypted_data_buf[670];   // modexp_top.v(222)
    assign encrypted_data_buf_next[669] = exp_valid ? exp_out[669] : encrypted_data_buf[669];   // modexp_top.v(222)
    assign encrypted_data_buf_next[668] = exp_valid ? exp_out[668] : encrypted_data_buf[668];   // modexp_top.v(222)
    assign encrypted_data_buf_next[667] = exp_valid ? exp_out[667] : encrypted_data_buf[667];   // modexp_top.v(222)
    assign encrypted_data_buf_next[666] = exp_valid ? exp_out[666] : encrypted_data_buf[666];   // modexp_top.v(222)
    assign encrypted_data_buf_next[665] = exp_valid ? exp_out[665] : encrypted_data_buf[665];   // modexp_top.v(222)
    assign encrypted_data_buf_next[664] = exp_valid ? exp_out[664] : encrypted_data_buf[664];   // modexp_top.v(222)
    assign encrypted_data_buf_next[663] = exp_valid ? exp_out[663] : encrypted_data_buf[663];   // modexp_top.v(222)
    assign encrypted_data_buf_next[662] = exp_valid ? exp_out[662] : encrypted_data_buf[662];   // modexp_top.v(222)
    assign encrypted_data_buf_next[661] = exp_valid ? exp_out[661] : encrypted_data_buf[661];   // modexp_top.v(222)
    assign encrypted_data_buf_next[660] = exp_valid ? exp_out[660] : encrypted_data_buf[660];   // modexp_top.v(222)
    assign encrypted_data_buf_next[659] = exp_valid ? exp_out[659] : encrypted_data_buf[659];   // modexp_top.v(222)
    assign encrypted_data_buf_next[658] = exp_valid ? exp_out[658] : encrypted_data_buf[658];   // modexp_top.v(222)
    assign encrypted_data_buf_next[657] = exp_valid ? exp_out[657] : encrypted_data_buf[657];   // modexp_top.v(222)
    assign encrypted_data_buf_next[656] = exp_valid ? exp_out[656] : encrypted_data_buf[656];   // modexp_top.v(222)
    assign encrypted_data_buf_next[655] = exp_valid ? exp_out[655] : encrypted_data_buf[655];   // modexp_top.v(222)
    assign encrypted_data_buf_next[654] = exp_valid ? exp_out[654] : encrypted_data_buf[654];   // modexp_top.v(222)
    assign encrypted_data_buf_next[653] = exp_valid ? exp_out[653] : encrypted_data_buf[653];   // modexp_top.v(222)
    assign encrypted_data_buf_next[652] = exp_valid ? exp_out[652] : encrypted_data_buf[652];   // modexp_top.v(222)
    assign encrypted_data_buf_next[651] = exp_valid ? exp_out[651] : encrypted_data_buf[651];   // modexp_top.v(222)
    assign encrypted_data_buf_next[650] = exp_valid ? exp_out[650] : encrypted_data_buf[650];   // modexp_top.v(222)
    assign encrypted_data_buf_next[649] = exp_valid ? exp_out[649] : encrypted_data_buf[649];   // modexp_top.v(222)
    assign encrypted_data_buf_next[648] = exp_valid ? exp_out[648] : encrypted_data_buf[648];   // modexp_top.v(222)
    assign encrypted_data_buf_next[647] = exp_valid ? exp_out[647] : encrypted_data_buf[647];   // modexp_top.v(222)
    assign encrypted_data_buf_next[646] = exp_valid ? exp_out[646] : encrypted_data_buf[646];   // modexp_top.v(222)
    assign encrypted_data_buf_next[645] = exp_valid ? exp_out[645] : encrypted_data_buf[645];   // modexp_top.v(222)
    assign encrypted_data_buf_next[644] = exp_valid ? exp_out[644] : encrypted_data_buf[644];   // modexp_top.v(222)
    assign encrypted_data_buf_next[643] = exp_valid ? exp_out[643] : encrypted_data_buf[643];   // modexp_top.v(222)
    assign encrypted_data_buf_next[642] = exp_valid ? exp_out[642] : encrypted_data_buf[642];   // modexp_top.v(222)
    assign encrypted_data_buf_next[641] = exp_valid ? exp_out[641] : encrypted_data_buf[641];   // modexp_top.v(222)
    assign encrypted_data_buf_next[640] = exp_valid ? exp_out[640] : encrypted_data_buf[640];   // modexp_top.v(222)
    assign encrypted_data_buf_next[639] = exp_valid ? exp_out[639] : encrypted_data_buf[639];   // modexp_top.v(222)
    assign encrypted_data_buf_next[638] = exp_valid ? exp_out[638] : encrypted_data_buf[638];   // modexp_top.v(222)
    assign encrypted_data_buf_next[637] = exp_valid ? exp_out[637] : encrypted_data_buf[637];   // modexp_top.v(222)
    assign encrypted_data_buf_next[636] = exp_valid ? exp_out[636] : encrypted_data_buf[636];   // modexp_top.v(222)
    assign encrypted_data_buf_next[635] = exp_valid ? exp_out[635] : encrypted_data_buf[635];   // modexp_top.v(222)
    assign encrypted_data_buf_next[634] = exp_valid ? exp_out[634] : encrypted_data_buf[634];   // modexp_top.v(222)
    assign encrypted_data_buf_next[633] = exp_valid ? exp_out[633] : encrypted_data_buf[633];   // modexp_top.v(222)
    assign encrypted_data_buf_next[632] = exp_valid ? exp_out[632] : encrypted_data_buf[632];   // modexp_top.v(222)
    assign encrypted_data_buf_next[631] = exp_valid ? exp_out[631] : encrypted_data_buf[631];   // modexp_top.v(222)
    assign encrypted_data_buf_next[630] = exp_valid ? exp_out[630] : encrypted_data_buf[630];   // modexp_top.v(222)
    assign encrypted_data_buf_next[629] = exp_valid ? exp_out[629] : encrypted_data_buf[629];   // modexp_top.v(222)
    assign encrypted_data_buf_next[628] = exp_valid ? exp_out[628] : encrypted_data_buf[628];   // modexp_top.v(222)
    assign encrypted_data_buf_next[627] = exp_valid ? exp_out[627] : encrypted_data_buf[627];   // modexp_top.v(222)
    assign encrypted_data_buf_next[626] = exp_valid ? exp_out[626] : encrypted_data_buf[626];   // modexp_top.v(222)
    assign encrypted_data_buf_next[625] = exp_valid ? exp_out[625] : encrypted_data_buf[625];   // modexp_top.v(222)
    assign encrypted_data_buf_next[624] = exp_valid ? exp_out[624] : encrypted_data_buf[624];   // modexp_top.v(222)
    assign encrypted_data_buf_next[623] = exp_valid ? exp_out[623] : encrypted_data_buf[623];   // modexp_top.v(222)
    assign encrypted_data_buf_next[622] = exp_valid ? exp_out[622] : encrypted_data_buf[622];   // modexp_top.v(222)
    assign encrypted_data_buf_next[621] = exp_valid ? exp_out[621] : encrypted_data_buf[621];   // modexp_top.v(222)
    assign encrypted_data_buf_next[620] = exp_valid ? exp_out[620] : encrypted_data_buf[620];   // modexp_top.v(222)
    assign encrypted_data_buf_next[619] = exp_valid ? exp_out[619] : encrypted_data_buf[619];   // modexp_top.v(222)
    assign encrypted_data_buf_next[618] = exp_valid ? exp_out[618] : encrypted_data_buf[618];   // modexp_top.v(222)
    assign encrypted_data_buf_next[617] = exp_valid ? exp_out[617] : encrypted_data_buf[617];   // modexp_top.v(222)
    assign encrypted_data_buf_next[616] = exp_valid ? exp_out[616] : encrypted_data_buf[616];   // modexp_top.v(222)
    assign encrypted_data_buf_next[615] = exp_valid ? exp_out[615] : encrypted_data_buf[615];   // modexp_top.v(222)
    assign encrypted_data_buf_next[614] = exp_valid ? exp_out[614] : encrypted_data_buf[614];   // modexp_top.v(222)
    assign encrypted_data_buf_next[613] = exp_valid ? exp_out[613] : encrypted_data_buf[613];   // modexp_top.v(222)
    assign encrypted_data_buf_next[612] = exp_valid ? exp_out[612] : encrypted_data_buf[612];   // modexp_top.v(222)
    assign encrypted_data_buf_next[611] = exp_valid ? exp_out[611] : encrypted_data_buf[611];   // modexp_top.v(222)
    assign encrypted_data_buf_next[610] = exp_valid ? exp_out[610] : encrypted_data_buf[610];   // modexp_top.v(222)
    assign encrypted_data_buf_next[609] = exp_valid ? exp_out[609] : encrypted_data_buf[609];   // modexp_top.v(222)
    assign encrypted_data_buf_next[608] = exp_valid ? exp_out[608] : encrypted_data_buf[608];   // modexp_top.v(222)
    assign encrypted_data_buf_next[607] = exp_valid ? exp_out[607] : encrypted_data_buf[607];   // modexp_top.v(222)
    assign encrypted_data_buf_next[606] = exp_valid ? exp_out[606] : encrypted_data_buf[606];   // modexp_top.v(222)
    assign encrypted_data_buf_next[605] = exp_valid ? exp_out[605] : encrypted_data_buf[605];   // modexp_top.v(222)
    assign encrypted_data_buf_next[604] = exp_valid ? exp_out[604] : encrypted_data_buf[604];   // modexp_top.v(222)
    assign encrypted_data_buf_next[603] = exp_valid ? exp_out[603] : encrypted_data_buf[603];   // modexp_top.v(222)
    assign encrypted_data_buf_next[602] = exp_valid ? exp_out[602] : encrypted_data_buf[602];   // modexp_top.v(222)
    assign encrypted_data_buf_next[601] = exp_valid ? exp_out[601] : encrypted_data_buf[601];   // modexp_top.v(222)
    assign encrypted_data_buf_next[600] = exp_valid ? exp_out[600] : encrypted_data_buf[600];   // modexp_top.v(222)
    assign encrypted_data_buf_next[599] = exp_valid ? exp_out[599] : encrypted_data_buf[599];   // modexp_top.v(222)
    assign encrypted_data_buf_next[598] = exp_valid ? exp_out[598] : encrypted_data_buf[598];   // modexp_top.v(222)
    assign encrypted_data_buf_next[597] = exp_valid ? exp_out[597] : encrypted_data_buf[597];   // modexp_top.v(222)
    assign encrypted_data_buf_next[596] = exp_valid ? exp_out[596] : encrypted_data_buf[596];   // modexp_top.v(222)
    assign encrypted_data_buf_next[595] = exp_valid ? exp_out[595] : encrypted_data_buf[595];   // modexp_top.v(222)
    assign encrypted_data_buf_next[594] = exp_valid ? exp_out[594] : encrypted_data_buf[594];   // modexp_top.v(222)
    assign encrypted_data_buf_next[593] = exp_valid ? exp_out[593] : encrypted_data_buf[593];   // modexp_top.v(222)
    assign encrypted_data_buf_next[592] = exp_valid ? exp_out[592] : encrypted_data_buf[592];   // modexp_top.v(222)
    assign encrypted_data_buf_next[591] = exp_valid ? exp_out[591] : encrypted_data_buf[591];   // modexp_top.v(222)
    assign encrypted_data_buf_next[590] = exp_valid ? exp_out[590] : encrypted_data_buf[590];   // modexp_top.v(222)
    assign encrypted_data_buf_next[589] = exp_valid ? exp_out[589] : encrypted_data_buf[589];   // modexp_top.v(222)
    assign encrypted_data_buf_next[588] = exp_valid ? exp_out[588] : encrypted_data_buf[588];   // modexp_top.v(222)
    assign encrypted_data_buf_next[587] = exp_valid ? exp_out[587] : encrypted_data_buf[587];   // modexp_top.v(222)
    assign encrypted_data_buf_next[586] = exp_valid ? exp_out[586] : encrypted_data_buf[586];   // modexp_top.v(222)
    assign encrypted_data_buf_next[585] = exp_valid ? exp_out[585] : encrypted_data_buf[585];   // modexp_top.v(222)
    assign encrypted_data_buf_next[584] = exp_valid ? exp_out[584] : encrypted_data_buf[584];   // modexp_top.v(222)
    assign encrypted_data_buf_next[583] = exp_valid ? exp_out[583] : encrypted_data_buf[583];   // modexp_top.v(222)
    assign encrypted_data_buf_next[582] = exp_valid ? exp_out[582] : encrypted_data_buf[582];   // modexp_top.v(222)
    assign encrypted_data_buf_next[581] = exp_valid ? exp_out[581] : encrypted_data_buf[581];   // modexp_top.v(222)
    assign encrypted_data_buf_next[580] = exp_valid ? exp_out[580] : encrypted_data_buf[580];   // modexp_top.v(222)
    assign encrypted_data_buf_next[579] = exp_valid ? exp_out[579] : encrypted_data_buf[579];   // modexp_top.v(222)
    assign encrypted_data_buf_next[578] = exp_valid ? exp_out[578] : encrypted_data_buf[578];   // modexp_top.v(222)
    assign encrypted_data_buf_next[577] = exp_valid ? exp_out[577] : encrypted_data_buf[577];   // modexp_top.v(222)
    assign encrypted_data_buf_next[576] = exp_valid ? exp_out[576] : encrypted_data_buf[576];   // modexp_top.v(222)
    assign encrypted_data_buf_next[575] = exp_valid ? exp_out[575] : encrypted_data_buf[575];   // modexp_top.v(222)
    assign encrypted_data_buf_next[574] = exp_valid ? exp_out[574] : encrypted_data_buf[574];   // modexp_top.v(222)
    assign encrypted_data_buf_next[573] = exp_valid ? exp_out[573] : encrypted_data_buf[573];   // modexp_top.v(222)
    assign encrypted_data_buf_next[572] = exp_valid ? exp_out[572] : encrypted_data_buf[572];   // modexp_top.v(222)
    assign encrypted_data_buf_next[571] = exp_valid ? exp_out[571] : encrypted_data_buf[571];   // modexp_top.v(222)
    assign encrypted_data_buf_next[570] = exp_valid ? exp_out[570] : encrypted_data_buf[570];   // modexp_top.v(222)
    assign encrypted_data_buf_next[569] = exp_valid ? exp_out[569] : encrypted_data_buf[569];   // modexp_top.v(222)
    assign encrypted_data_buf_next[568] = exp_valid ? exp_out[568] : encrypted_data_buf[568];   // modexp_top.v(222)
    assign encrypted_data_buf_next[567] = exp_valid ? exp_out[567] : encrypted_data_buf[567];   // modexp_top.v(222)
    assign encrypted_data_buf_next[566] = exp_valid ? exp_out[566] : encrypted_data_buf[566];   // modexp_top.v(222)
    assign encrypted_data_buf_next[565] = exp_valid ? exp_out[565] : encrypted_data_buf[565];   // modexp_top.v(222)
    assign encrypted_data_buf_next[564] = exp_valid ? exp_out[564] : encrypted_data_buf[564];   // modexp_top.v(222)
    assign encrypted_data_buf_next[563] = exp_valid ? exp_out[563] : encrypted_data_buf[563];   // modexp_top.v(222)
    assign encrypted_data_buf_next[562] = exp_valid ? exp_out[562] : encrypted_data_buf[562];   // modexp_top.v(222)
    assign encrypted_data_buf_next[561] = exp_valid ? exp_out[561] : encrypted_data_buf[561];   // modexp_top.v(222)
    assign encrypted_data_buf_next[560] = exp_valid ? exp_out[560] : encrypted_data_buf[560];   // modexp_top.v(222)
    assign encrypted_data_buf_next[559] = exp_valid ? exp_out[559] : encrypted_data_buf[559];   // modexp_top.v(222)
    assign encrypted_data_buf_next[558] = exp_valid ? exp_out[558] : encrypted_data_buf[558];   // modexp_top.v(222)
    assign encrypted_data_buf_next[557] = exp_valid ? exp_out[557] : encrypted_data_buf[557];   // modexp_top.v(222)
    assign encrypted_data_buf_next[556] = exp_valid ? exp_out[556] : encrypted_data_buf[556];   // modexp_top.v(222)
    assign encrypted_data_buf_next[555] = exp_valid ? exp_out[555] : encrypted_data_buf[555];   // modexp_top.v(222)
    assign encrypted_data_buf_next[554] = exp_valid ? exp_out[554] : encrypted_data_buf[554];   // modexp_top.v(222)
    assign encrypted_data_buf_next[553] = exp_valid ? exp_out[553] : encrypted_data_buf[553];   // modexp_top.v(222)
    assign encrypted_data_buf_next[552] = exp_valid ? exp_out[552] : encrypted_data_buf[552];   // modexp_top.v(222)
    assign encrypted_data_buf_next[551] = exp_valid ? exp_out[551] : encrypted_data_buf[551];   // modexp_top.v(222)
    assign encrypted_data_buf_next[550] = exp_valid ? exp_out[550] : encrypted_data_buf[550];   // modexp_top.v(222)
    assign encrypted_data_buf_next[549] = exp_valid ? exp_out[549] : encrypted_data_buf[549];   // modexp_top.v(222)
    assign encrypted_data_buf_next[548] = exp_valid ? exp_out[548] : encrypted_data_buf[548];   // modexp_top.v(222)
    assign encrypted_data_buf_next[547] = exp_valid ? exp_out[547] : encrypted_data_buf[547];   // modexp_top.v(222)
    assign encrypted_data_buf_next[546] = exp_valid ? exp_out[546] : encrypted_data_buf[546];   // modexp_top.v(222)
    assign encrypted_data_buf_next[545] = exp_valid ? exp_out[545] : encrypted_data_buf[545];   // modexp_top.v(222)
    assign encrypted_data_buf_next[544] = exp_valid ? exp_out[544] : encrypted_data_buf[544];   // modexp_top.v(222)
    assign encrypted_data_buf_next[543] = exp_valid ? exp_out[543] : encrypted_data_buf[543];   // modexp_top.v(222)
    assign encrypted_data_buf_next[542] = exp_valid ? exp_out[542] : encrypted_data_buf[542];   // modexp_top.v(222)
    assign encrypted_data_buf_next[541] = exp_valid ? exp_out[541] : encrypted_data_buf[541];   // modexp_top.v(222)
    assign encrypted_data_buf_next[540] = exp_valid ? exp_out[540] : encrypted_data_buf[540];   // modexp_top.v(222)
    assign encrypted_data_buf_next[539] = exp_valid ? exp_out[539] : encrypted_data_buf[539];   // modexp_top.v(222)
    assign encrypted_data_buf_next[538] = exp_valid ? exp_out[538] : encrypted_data_buf[538];   // modexp_top.v(222)
    assign encrypted_data_buf_next[537] = exp_valid ? exp_out[537] : encrypted_data_buf[537];   // modexp_top.v(222)
    assign encrypted_data_buf_next[536] = exp_valid ? exp_out[536] : encrypted_data_buf[536];   // modexp_top.v(222)
    assign encrypted_data_buf_next[535] = exp_valid ? exp_out[535] : encrypted_data_buf[535];   // modexp_top.v(222)
    assign encrypted_data_buf_next[534] = exp_valid ? exp_out[534] : encrypted_data_buf[534];   // modexp_top.v(222)
    assign encrypted_data_buf_next[533] = exp_valid ? exp_out[533] : encrypted_data_buf[533];   // modexp_top.v(222)
    assign encrypted_data_buf_next[532] = exp_valid ? exp_out[532] : encrypted_data_buf[532];   // modexp_top.v(222)
    assign encrypted_data_buf_next[531] = exp_valid ? exp_out[531] : encrypted_data_buf[531];   // modexp_top.v(222)
    assign encrypted_data_buf_next[530] = exp_valid ? exp_out[530] : encrypted_data_buf[530];   // modexp_top.v(222)
    assign encrypted_data_buf_next[529] = exp_valid ? exp_out[529] : encrypted_data_buf[529];   // modexp_top.v(222)
    assign encrypted_data_buf_next[528] = exp_valid ? exp_out[528] : encrypted_data_buf[528];   // modexp_top.v(222)
    assign encrypted_data_buf_next[527] = exp_valid ? exp_out[527] : encrypted_data_buf[527];   // modexp_top.v(222)
    assign encrypted_data_buf_next[526] = exp_valid ? exp_out[526] : encrypted_data_buf[526];   // modexp_top.v(222)
    assign encrypted_data_buf_next[525] = exp_valid ? exp_out[525] : encrypted_data_buf[525];   // modexp_top.v(222)
    assign encrypted_data_buf_next[524] = exp_valid ? exp_out[524] : encrypted_data_buf[524];   // modexp_top.v(222)
    assign encrypted_data_buf_next[523] = exp_valid ? exp_out[523] : encrypted_data_buf[523];   // modexp_top.v(222)
    assign encrypted_data_buf_next[522] = exp_valid ? exp_out[522] : encrypted_data_buf[522];   // modexp_top.v(222)
    assign encrypted_data_buf_next[521] = exp_valid ? exp_out[521] : encrypted_data_buf[521];   // modexp_top.v(222)
    assign encrypted_data_buf_next[520] = exp_valid ? exp_out[520] : encrypted_data_buf[520];   // modexp_top.v(222)
    assign encrypted_data_buf_next[519] = exp_valid ? exp_out[519] : encrypted_data_buf[519];   // modexp_top.v(222)
    assign encrypted_data_buf_next[518] = exp_valid ? exp_out[518] : encrypted_data_buf[518];   // modexp_top.v(222)
    assign encrypted_data_buf_next[517] = exp_valid ? exp_out[517] : encrypted_data_buf[517];   // modexp_top.v(222)
    assign encrypted_data_buf_next[516] = exp_valid ? exp_out[516] : encrypted_data_buf[516];   // modexp_top.v(222)
    assign encrypted_data_buf_next[515] = exp_valid ? exp_out[515] : encrypted_data_buf[515];   // modexp_top.v(222)
    assign encrypted_data_buf_next[514] = exp_valid ? exp_out[514] : encrypted_data_buf[514];   // modexp_top.v(222)
    assign encrypted_data_buf_next[513] = exp_valid ? exp_out[513] : encrypted_data_buf[513];   // modexp_top.v(222)
    assign encrypted_data_buf_next[512] = exp_valid ? exp_out[512] : encrypted_data_buf[512];   // modexp_top.v(222)
    assign encrypted_data_buf_next[511] = exp_valid ? exp_out[511] : encrypted_data_buf[511];   // modexp_top.v(222)
    assign encrypted_data_buf_next[510] = exp_valid ? exp_out[510] : encrypted_data_buf[510];   // modexp_top.v(222)
    assign encrypted_data_buf_next[509] = exp_valid ? exp_out[509] : encrypted_data_buf[509];   // modexp_top.v(222)
    assign encrypted_data_buf_next[508] = exp_valid ? exp_out[508] : encrypted_data_buf[508];   // modexp_top.v(222)
    assign encrypted_data_buf_next[507] = exp_valid ? exp_out[507] : encrypted_data_buf[507];   // modexp_top.v(222)
    assign encrypted_data_buf_next[506] = exp_valid ? exp_out[506] : encrypted_data_buf[506];   // modexp_top.v(222)
    assign encrypted_data_buf_next[505] = exp_valid ? exp_out[505] : encrypted_data_buf[505];   // modexp_top.v(222)
    assign encrypted_data_buf_next[504] = exp_valid ? exp_out[504] : encrypted_data_buf[504];   // modexp_top.v(222)
    assign encrypted_data_buf_next[503] = exp_valid ? exp_out[503] : encrypted_data_buf[503];   // modexp_top.v(222)
    assign encrypted_data_buf_next[502] = exp_valid ? exp_out[502] : encrypted_data_buf[502];   // modexp_top.v(222)
    assign encrypted_data_buf_next[501] = exp_valid ? exp_out[501] : encrypted_data_buf[501];   // modexp_top.v(222)
    assign encrypted_data_buf_next[500] = exp_valid ? exp_out[500] : encrypted_data_buf[500];   // modexp_top.v(222)
    assign encrypted_data_buf_next[499] = exp_valid ? exp_out[499] : encrypted_data_buf[499];   // modexp_top.v(222)
    assign encrypted_data_buf_next[498] = exp_valid ? exp_out[498] : encrypted_data_buf[498];   // modexp_top.v(222)
    assign encrypted_data_buf_next[497] = exp_valid ? exp_out[497] : encrypted_data_buf[497];   // modexp_top.v(222)
    assign encrypted_data_buf_next[496] = exp_valid ? exp_out[496] : encrypted_data_buf[496];   // modexp_top.v(222)
    assign encrypted_data_buf_next[495] = exp_valid ? exp_out[495] : encrypted_data_buf[495];   // modexp_top.v(222)
    assign encrypted_data_buf_next[494] = exp_valid ? exp_out[494] : encrypted_data_buf[494];   // modexp_top.v(222)
    assign encrypted_data_buf_next[493] = exp_valid ? exp_out[493] : encrypted_data_buf[493];   // modexp_top.v(222)
    assign encrypted_data_buf_next[492] = exp_valid ? exp_out[492] : encrypted_data_buf[492];   // modexp_top.v(222)
    assign encrypted_data_buf_next[491] = exp_valid ? exp_out[491] : encrypted_data_buf[491];   // modexp_top.v(222)
    assign encrypted_data_buf_next[490] = exp_valid ? exp_out[490] : encrypted_data_buf[490];   // modexp_top.v(222)
    assign encrypted_data_buf_next[489] = exp_valid ? exp_out[489] : encrypted_data_buf[489];   // modexp_top.v(222)
    assign encrypted_data_buf_next[488] = exp_valid ? exp_out[488] : encrypted_data_buf[488];   // modexp_top.v(222)
    assign encrypted_data_buf_next[487] = exp_valid ? exp_out[487] : encrypted_data_buf[487];   // modexp_top.v(222)
    assign encrypted_data_buf_next[486] = exp_valid ? exp_out[486] : encrypted_data_buf[486];   // modexp_top.v(222)
    assign encrypted_data_buf_next[485] = exp_valid ? exp_out[485] : encrypted_data_buf[485];   // modexp_top.v(222)
    assign encrypted_data_buf_next[484] = exp_valid ? exp_out[484] : encrypted_data_buf[484];   // modexp_top.v(222)
    assign encrypted_data_buf_next[483] = exp_valid ? exp_out[483] : encrypted_data_buf[483];   // modexp_top.v(222)
    assign encrypted_data_buf_next[482] = exp_valid ? exp_out[482] : encrypted_data_buf[482];   // modexp_top.v(222)
    assign encrypted_data_buf_next[481] = exp_valid ? exp_out[481] : encrypted_data_buf[481];   // modexp_top.v(222)
    assign encrypted_data_buf_next[480] = exp_valid ? exp_out[480] : encrypted_data_buf[480];   // modexp_top.v(222)
    assign encrypted_data_buf_next[479] = exp_valid ? exp_out[479] : encrypted_data_buf[479];   // modexp_top.v(222)
    assign encrypted_data_buf_next[478] = exp_valid ? exp_out[478] : encrypted_data_buf[478];   // modexp_top.v(222)
    assign encrypted_data_buf_next[477] = exp_valid ? exp_out[477] : encrypted_data_buf[477];   // modexp_top.v(222)
    assign encrypted_data_buf_next[476] = exp_valid ? exp_out[476] : encrypted_data_buf[476];   // modexp_top.v(222)
    assign encrypted_data_buf_next[475] = exp_valid ? exp_out[475] : encrypted_data_buf[475];   // modexp_top.v(222)
    assign encrypted_data_buf_next[474] = exp_valid ? exp_out[474] : encrypted_data_buf[474];   // modexp_top.v(222)
    assign encrypted_data_buf_next[473] = exp_valid ? exp_out[473] : encrypted_data_buf[473];   // modexp_top.v(222)
    assign encrypted_data_buf_next[472] = exp_valid ? exp_out[472] : encrypted_data_buf[472];   // modexp_top.v(222)
    assign encrypted_data_buf_next[471] = exp_valid ? exp_out[471] : encrypted_data_buf[471];   // modexp_top.v(222)
    assign encrypted_data_buf_next[470] = exp_valid ? exp_out[470] : encrypted_data_buf[470];   // modexp_top.v(222)
    assign encrypted_data_buf_next[469] = exp_valid ? exp_out[469] : encrypted_data_buf[469];   // modexp_top.v(222)
    assign encrypted_data_buf_next[468] = exp_valid ? exp_out[468] : encrypted_data_buf[468];   // modexp_top.v(222)
    assign encrypted_data_buf_next[467] = exp_valid ? exp_out[467] : encrypted_data_buf[467];   // modexp_top.v(222)
    assign encrypted_data_buf_next[466] = exp_valid ? exp_out[466] : encrypted_data_buf[466];   // modexp_top.v(222)
    assign encrypted_data_buf_next[465] = exp_valid ? exp_out[465] : encrypted_data_buf[465];   // modexp_top.v(222)
    assign encrypted_data_buf_next[464] = exp_valid ? exp_out[464] : encrypted_data_buf[464];   // modexp_top.v(222)
    assign encrypted_data_buf_next[463] = exp_valid ? exp_out[463] : encrypted_data_buf[463];   // modexp_top.v(222)
    assign encrypted_data_buf_next[462] = exp_valid ? exp_out[462] : encrypted_data_buf[462];   // modexp_top.v(222)
    assign encrypted_data_buf_next[461] = exp_valid ? exp_out[461] : encrypted_data_buf[461];   // modexp_top.v(222)
    assign encrypted_data_buf_next[460] = exp_valid ? exp_out[460] : encrypted_data_buf[460];   // modexp_top.v(222)
    assign encrypted_data_buf_next[459] = exp_valid ? exp_out[459] : encrypted_data_buf[459];   // modexp_top.v(222)
    assign encrypted_data_buf_next[458] = exp_valid ? exp_out[458] : encrypted_data_buf[458];   // modexp_top.v(222)
    assign encrypted_data_buf_next[457] = exp_valid ? exp_out[457] : encrypted_data_buf[457];   // modexp_top.v(222)
    assign encrypted_data_buf_next[456] = exp_valid ? exp_out[456] : encrypted_data_buf[456];   // modexp_top.v(222)
    assign encrypted_data_buf_next[455] = exp_valid ? exp_out[455] : encrypted_data_buf[455];   // modexp_top.v(222)
    assign encrypted_data_buf_next[454] = exp_valid ? exp_out[454] : encrypted_data_buf[454];   // modexp_top.v(222)
    assign encrypted_data_buf_next[453] = exp_valid ? exp_out[453] : encrypted_data_buf[453];   // modexp_top.v(222)
    assign encrypted_data_buf_next[452] = exp_valid ? exp_out[452] : encrypted_data_buf[452];   // modexp_top.v(222)
    assign encrypted_data_buf_next[451] = exp_valid ? exp_out[451] : encrypted_data_buf[451];   // modexp_top.v(222)
    assign encrypted_data_buf_next[450] = exp_valid ? exp_out[450] : encrypted_data_buf[450];   // modexp_top.v(222)
    assign encrypted_data_buf_next[449] = exp_valid ? exp_out[449] : encrypted_data_buf[449];   // modexp_top.v(222)
    assign encrypted_data_buf_next[448] = exp_valid ? exp_out[448] : encrypted_data_buf[448];   // modexp_top.v(222)
    assign encrypted_data_buf_next[447] = exp_valid ? exp_out[447] : encrypted_data_buf[447];   // modexp_top.v(222)
    assign encrypted_data_buf_next[446] = exp_valid ? exp_out[446] : encrypted_data_buf[446];   // modexp_top.v(222)
    assign encrypted_data_buf_next[445] = exp_valid ? exp_out[445] : encrypted_data_buf[445];   // modexp_top.v(222)
    assign encrypted_data_buf_next[444] = exp_valid ? exp_out[444] : encrypted_data_buf[444];   // modexp_top.v(222)
    assign encrypted_data_buf_next[443] = exp_valid ? exp_out[443] : encrypted_data_buf[443];   // modexp_top.v(222)
    assign encrypted_data_buf_next[442] = exp_valid ? exp_out[442] : encrypted_data_buf[442];   // modexp_top.v(222)
    assign encrypted_data_buf_next[441] = exp_valid ? exp_out[441] : encrypted_data_buf[441];   // modexp_top.v(222)
    assign encrypted_data_buf_next[440] = exp_valid ? exp_out[440] : encrypted_data_buf[440];   // modexp_top.v(222)
    assign encrypted_data_buf_next[439] = exp_valid ? exp_out[439] : encrypted_data_buf[439];   // modexp_top.v(222)
    assign encrypted_data_buf_next[438] = exp_valid ? exp_out[438] : encrypted_data_buf[438];   // modexp_top.v(222)
    assign encrypted_data_buf_next[437] = exp_valid ? exp_out[437] : encrypted_data_buf[437];   // modexp_top.v(222)
    assign encrypted_data_buf_next[436] = exp_valid ? exp_out[436] : encrypted_data_buf[436];   // modexp_top.v(222)
    assign encrypted_data_buf_next[435] = exp_valid ? exp_out[435] : encrypted_data_buf[435];   // modexp_top.v(222)
    assign encrypted_data_buf_next[434] = exp_valid ? exp_out[434] : encrypted_data_buf[434];   // modexp_top.v(222)
    assign encrypted_data_buf_next[433] = exp_valid ? exp_out[433] : encrypted_data_buf[433];   // modexp_top.v(222)
    assign encrypted_data_buf_next[432] = exp_valid ? exp_out[432] : encrypted_data_buf[432];   // modexp_top.v(222)
    assign encrypted_data_buf_next[431] = exp_valid ? exp_out[431] : encrypted_data_buf[431];   // modexp_top.v(222)
    assign encrypted_data_buf_next[430] = exp_valid ? exp_out[430] : encrypted_data_buf[430];   // modexp_top.v(222)
    assign encrypted_data_buf_next[429] = exp_valid ? exp_out[429] : encrypted_data_buf[429];   // modexp_top.v(222)
    assign encrypted_data_buf_next[428] = exp_valid ? exp_out[428] : encrypted_data_buf[428];   // modexp_top.v(222)
    assign encrypted_data_buf_next[427] = exp_valid ? exp_out[427] : encrypted_data_buf[427];   // modexp_top.v(222)
    assign encrypted_data_buf_next[426] = exp_valid ? exp_out[426] : encrypted_data_buf[426];   // modexp_top.v(222)
    assign encrypted_data_buf_next[425] = exp_valid ? exp_out[425] : encrypted_data_buf[425];   // modexp_top.v(222)
    assign encrypted_data_buf_next[424] = exp_valid ? exp_out[424] : encrypted_data_buf[424];   // modexp_top.v(222)
    assign encrypted_data_buf_next[423] = exp_valid ? exp_out[423] : encrypted_data_buf[423];   // modexp_top.v(222)
    assign encrypted_data_buf_next[422] = exp_valid ? exp_out[422] : encrypted_data_buf[422];   // modexp_top.v(222)
    assign encrypted_data_buf_next[421] = exp_valid ? exp_out[421] : encrypted_data_buf[421];   // modexp_top.v(222)
    assign encrypted_data_buf_next[420] = exp_valid ? exp_out[420] : encrypted_data_buf[420];   // modexp_top.v(222)
    assign encrypted_data_buf_next[419] = exp_valid ? exp_out[419] : encrypted_data_buf[419];   // modexp_top.v(222)
    assign encrypted_data_buf_next[418] = exp_valid ? exp_out[418] : encrypted_data_buf[418];   // modexp_top.v(222)
    assign encrypted_data_buf_next[417] = exp_valid ? exp_out[417] : encrypted_data_buf[417];   // modexp_top.v(222)
    assign encrypted_data_buf_next[416] = exp_valid ? exp_out[416] : encrypted_data_buf[416];   // modexp_top.v(222)
    assign encrypted_data_buf_next[415] = exp_valid ? exp_out[415] : encrypted_data_buf[415];   // modexp_top.v(222)
    assign encrypted_data_buf_next[414] = exp_valid ? exp_out[414] : encrypted_data_buf[414];   // modexp_top.v(222)
    assign encrypted_data_buf_next[413] = exp_valid ? exp_out[413] : encrypted_data_buf[413];   // modexp_top.v(222)
    assign encrypted_data_buf_next[412] = exp_valid ? exp_out[412] : encrypted_data_buf[412];   // modexp_top.v(222)
    assign encrypted_data_buf_next[411] = exp_valid ? exp_out[411] : encrypted_data_buf[411];   // modexp_top.v(222)
    assign encrypted_data_buf_next[410] = exp_valid ? exp_out[410] : encrypted_data_buf[410];   // modexp_top.v(222)
    assign encrypted_data_buf_next[409] = exp_valid ? exp_out[409] : encrypted_data_buf[409];   // modexp_top.v(222)
    assign encrypted_data_buf_next[408] = exp_valid ? exp_out[408] : encrypted_data_buf[408];   // modexp_top.v(222)
    assign encrypted_data_buf_next[407] = exp_valid ? exp_out[407] : encrypted_data_buf[407];   // modexp_top.v(222)
    assign encrypted_data_buf_next[406] = exp_valid ? exp_out[406] : encrypted_data_buf[406];   // modexp_top.v(222)
    assign encrypted_data_buf_next[405] = exp_valid ? exp_out[405] : encrypted_data_buf[405];   // modexp_top.v(222)
    assign encrypted_data_buf_next[404] = exp_valid ? exp_out[404] : encrypted_data_buf[404];   // modexp_top.v(222)
    assign encrypted_data_buf_next[403] = exp_valid ? exp_out[403] : encrypted_data_buf[403];   // modexp_top.v(222)
    assign encrypted_data_buf_next[402] = exp_valid ? exp_out[402] : encrypted_data_buf[402];   // modexp_top.v(222)
    assign encrypted_data_buf_next[401] = exp_valid ? exp_out[401] : encrypted_data_buf[401];   // modexp_top.v(222)
    assign encrypted_data_buf_next[400] = exp_valid ? exp_out[400] : encrypted_data_buf[400];   // modexp_top.v(222)
    assign encrypted_data_buf_next[399] = exp_valid ? exp_out[399] : encrypted_data_buf[399];   // modexp_top.v(222)
    assign encrypted_data_buf_next[398] = exp_valid ? exp_out[398] : encrypted_data_buf[398];   // modexp_top.v(222)
    assign encrypted_data_buf_next[397] = exp_valid ? exp_out[397] : encrypted_data_buf[397];   // modexp_top.v(222)
    assign encrypted_data_buf_next[396] = exp_valid ? exp_out[396] : encrypted_data_buf[396];   // modexp_top.v(222)
    assign encrypted_data_buf_next[395] = exp_valid ? exp_out[395] : encrypted_data_buf[395];   // modexp_top.v(222)
    assign encrypted_data_buf_next[394] = exp_valid ? exp_out[394] : encrypted_data_buf[394];   // modexp_top.v(222)
    assign encrypted_data_buf_next[393] = exp_valid ? exp_out[393] : encrypted_data_buf[393];   // modexp_top.v(222)
    assign encrypted_data_buf_next[392] = exp_valid ? exp_out[392] : encrypted_data_buf[392];   // modexp_top.v(222)
    assign encrypted_data_buf_next[391] = exp_valid ? exp_out[391] : encrypted_data_buf[391];   // modexp_top.v(222)
    assign encrypted_data_buf_next[390] = exp_valid ? exp_out[390] : encrypted_data_buf[390];   // modexp_top.v(222)
    assign encrypted_data_buf_next[389] = exp_valid ? exp_out[389] : encrypted_data_buf[389];   // modexp_top.v(222)
    assign encrypted_data_buf_next[388] = exp_valid ? exp_out[388] : encrypted_data_buf[388];   // modexp_top.v(222)
    assign encrypted_data_buf_next[387] = exp_valid ? exp_out[387] : encrypted_data_buf[387];   // modexp_top.v(222)
    assign encrypted_data_buf_next[386] = exp_valid ? exp_out[386] : encrypted_data_buf[386];   // modexp_top.v(222)
    assign encrypted_data_buf_next[385] = exp_valid ? exp_out[385] : encrypted_data_buf[385];   // modexp_top.v(222)
    assign encrypted_data_buf_next[384] = exp_valid ? exp_out[384] : encrypted_data_buf[384];   // modexp_top.v(222)
    assign encrypted_data_buf_next[383] = exp_valid ? exp_out[383] : encrypted_data_buf[383];   // modexp_top.v(222)
    assign encrypted_data_buf_next[382] = exp_valid ? exp_out[382] : encrypted_data_buf[382];   // modexp_top.v(222)
    assign encrypted_data_buf_next[381] = exp_valid ? exp_out[381] : encrypted_data_buf[381];   // modexp_top.v(222)
    assign encrypted_data_buf_next[380] = exp_valid ? exp_out[380] : encrypted_data_buf[380];   // modexp_top.v(222)
    assign encrypted_data_buf_next[379] = exp_valid ? exp_out[379] : encrypted_data_buf[379];   // modexp_top.v(222)
    assign encrypted_data_buf_next[378] = exp_valid ? exp_out[378] : encrypted_data_buf[378];   // modexp_top.v(222)
    assign encrypted_data_buf_next[377] = exp_valid ? exp_out[377] : encrypted_data_buf[377];   // modexp_top.v(222)
    assign encrypted_data_buf_next[376] = exp_valid ? exp_out[376] : encrypted_data_buf[376];   // modexp_top.v(222)
    assign encrypted_data_buf_next[375] = exp_valid ? exp_out[375] : encrypted_data_buf[375];   // modexp_top.v(222)
    assign encrypted_data_buf_next[374] = exp_valid ? exp_out[374] : encrypted_data_buf[374];   // modexp_top.v(222)
    assign encrypted_data_buf_next[373] = exp_valid ? exp_out[373] : encrypted_data_buf[373];   // modexp_top.v(222)
    assign encrypted_data_buf_next[372] = exp_valid ? exp_out[372] : encrypted_data_buf[372];   // modexp_top.v(222)
    assign encrypted_data_buf_next[371] = exp_valid ? exp_out[371] : encrypted_data_buf[371];   // modexp_top.v(222)
    assign encrypted_data_buf_next[370] = exp_valid ? exp_out[370] : encrypted_data_buf[370];   // modexp_top.v(222)
    assign encrypted_data_buf_next[369] = exp_valid ? exp_out[369] : encrypted_data_buf[369];   // modexp_top.v(222)
    assign encrypted_data_buf_next[368] = exp_valid ? exp_out[368] : encrypted_data_buf[368];   // modexp_top.v(222)
    assign encrypted_data_buf_next[367] = exp_valid ? exp_out[367] : encrypted_data_buf[367];   // modexp_top.v(222)
    assign encrypted_data_buf_next[366] = exp_valid ? exp_out[366] : encrypted_data_buf[366];   // modexp_top.v(222)
    assign encrypted_data_buf_next[365] = exp_valid ? exp_out[365] : encrypted_data_buf[365];   // modexp_top.v(222)
    assign encrypted_data_buf_next[364] = exp_valid ? exp_out[364] : encrypted_data_buf[364];   // modexp_top.v(222)
    assign encrypted_data_buf_next[363] = exp_valid ? exp_out[363] : encrypted_data_buf[363];   // modexp_top.v(222)
    assign encrypted_data_buf_next[362] = exp_valid ? exp_out[362] : encrypted_data_buf[362];   // modexp_top.v(222)
    assign encrypted_data_buf_next[361] = exp_valid ? exp_out[361] : encrypted_data_buf[361];   // modexp_top.v(222)
    assign encrypted_data_buf_next[360] = exp_valid ? exp_out[360] : encrypted_data_buf[360];   // modexp_top.v(222)
    assign encrypted_data_buf_next[359] = exp_valid ? exp_out[359] : encrypted_data_buf[359];   // modexp_top.v(222)
    assign encrypted_data_buf_next[358] = exp_valid ? exp_out[358] : encrypted_data_buf[358];   // modexp_top.v(222)
    assign encrypted_data_buf_next[357] = exp_valid ? exp_out[357] : encrypted_data_buf[357];   // modexp_top.v(222)
    assign encrypted_data_buf_next[356] = exp_valid ? exp_out[356] : encrypted_data_buf[356];   // modexp_top.v(222)
    assign encrypted_data_buf_next[355] = exp_valid ? exp_out[355] : encrypted_data_buf[355];   // modexp_top.v(222)
    assign encrypted_data_buf_next[354] = exp_valid ? exp_out[354] : encrypted_data_buf[354];   // modexp_top.v(222)
    assign encrypted_data_buf_next[353] = exp_valid ? exp_out[353] : encrypted_data_buf[353];   // modexp_top.v(222)
    assign encrypted_data_buf_next[352] = exp_valid ? exp_out[352] : encrypted_data_buf[352];   // modexp_top.v(222)
    assign encrypted_data_buf_next[351] = exp_valid ? exp_out[351] : encrypted_data_buf[351];   // modexp_top.v(222)
    assign encrypted_data_buf_next[350] = exp_valid ? exp_out[350] : encrypted_data_buf[350];   // modexp_top.v(222)
    assign encrypted_data_buf_next[349] = exp_valid ? exp_out[349] : encrypted_data_buf[349];   // modexp_top.v(222)
    assign encrypted_data_buf_next[348] = exp_valid ? exp_out[348] : encrypted_data_buf[348];   // modexp_top.v(222)
    assign encrypted_data_buf_next[347] = exp_valid ? exp_out[347] : encrypted_data_buf[347];   // modexp_top.v(222)
    assign encrypted_data_buf_next[346] = exp_valid ? exp_out[346] : encrypted_data_buf[346];   // modexp_top.v(222)
    assign encrypted_data_buf_next[345] = exp_valid ? exp_out[345] : encrypted_data_buf[345];   // modexp_top.v(222)
    assign encrypted_data_buf_next[344] = exp_valid ? exp_out[344] : encrypted_data_buf[344];   // modexp_top.v(222)
    assign encrypted_data_buf_next[343] = exp_valid ? exp_out[343] : encrypted_data_buf[343];   // modexp_top.v(222)
    assign encrypted_data_buf_next[342] = exp_valid ? exp_out[342] : encrypted_data_buf[342];   // modexp_top.v(222)
    assign encrypted_data_buf_next[341] = exp_valid ? exp_out[341] : encrypted_data_buf[341];   // modexp_top.v(222)
    assign encrypted_data_buf_next[340] = exp_valid ? exp_out[340] : encrypted_data_buf[340];   // modexp_top.v(222)
    assign encrypted_data_buf_next[339] = exp_valid ? exp_out[339] : encrypted_data_buf[339];   // modexp_top.v(222)
    assign encrypted_data_buf_next[338] = exp_valid ? exp_out[338] : encrypted_data_buf[338];   // modexp_top.v(222)
    assign encrypted_data_buf_next[337] = exp_valid ? exp_out[337] : encrypted_data_buf[337];   // modexp_top.v(222)
    assign encrypted_data_buf_next[336] = exp_valid ? exp_out[336] : encrypted_data_buf[336];   // modexp_top.v(222)
    assign encrypted_data_buf_next[335] = exp_valid ? exp_out[335] : encrypted_data_buf[335];   // modexp_top.v(222)
    assign encrypted_data_buf_next[334] = exp_valid ? exp_out[334] : encrypted_data_buf[334];   // modexp_top.v(222)
    assign encrypted_data_buf_next[333] = exp_valid ? exp_out[333] : encrypted_data_buf[333];   // modexp_top.v(222)
    assign encrypted_data_buf_next[332] = exp_valid ? exp_out[332] : encrypted_data_buf[332];   // modexp_top.v(222)
    assign encrypted_data_buf_next[331] = exp_valid ? exp_out[331] : encrypted_data_buf[331];   // modexp_top.v(222)
    assign encrypted_data_buf_next[330] = exp_valid ? exp_out[330] : encrypted_data_buf[330];   // modexp_top.v(222)
    assign encrypted_data_buf_next[329] = exp_valid ? exp_out[329] : encrypted_data_buf[329];   // modexp_top.v(222)
    assign encrypted_data_buf_next[328] = exp_valid ? exp_out[328] : encrypted_data_buf[328];   // modexp_top.v(222)
    assign encrypted_data_buf_next[327] = exp_valid ? exp_out[327] : encrypted_data_buf[327];   // modexp_top.v(222)
    assign encrypted_data_buf_next[326] = exp_valid ? exp_out[326] : encrypted_data_buf[326];   // modexp_top.v(222)
    assign encrypted_data_buf_next[325] = exp_valid ? exp_out[325] : encrypted_data_buf[325];   // modexp_top.v(222)
    assign encrypted_data_buf_next[324] = exp_valid ? exp_out[324] : encrypted_data_buf[324];   // modexp_top.v(222)
    assign encrypted_data_buf_next[323] = exp_valid ? exp_out[323] : encrypted_data_buf[323];   // modexp_top.v(222)
    assign encrypted_data_buf_next[322] = exp_valid ? exp_out[322] : encrypted_data_buf[322];   // modexp_top.v(222)
    assign encrypted_data_buf_next[321] = exp_valid ? exp_out[321] : encrypted_data_buf[321];   // modexp_top.v(222)
    assign encrypted_data_buf_next[320] = exp_valid ? exp_out[320] : encrypted_data_buf[320];   // modexp_top.v(222)
    assign encrypted_data_buf_next[319] = exp_valid ? exp_out[319] : encrypted_data_buf[319];   // modexp_top.v(222)
    assign encrypted_data_buf_next[318] = exp_valid ? exp_out[318] : encrypted_data_buf[318];   // modexp_top.v(222)
    assign encrypted_data_buf_next[317] = exp_valid ? exp_out[317] : encrypted_data_buf[317];   // modexp_top.v(222)
    assign encrypted_data_buf_next[316] = exp_valid ? exp_out[316] : encrypted_data_buf[316];   // modexp_top.v(222)
    assign encrypted_data_buf_next[315] = exp_valid ? exp_out[315] : encrypted_data_buf[315];   // modexp_top.v(222)
    assign encrypted_data_buf_next[314] = exp_valid ? exp_out[314] : encrypted_data_buf[314];   // modexp_top.v(222)
    assign encrypted_data_buf_next[313] = exp_valid ? exp_out[313] : encrypted_data_buf[313];   // modexp_top.v(222)
    assign encrypted_data_buf_next[312] = exp_valid ? exp_out[312] : encrypted_data_buf[312];   // modexp_top.v(222)
    assign encrypted_data_buf_next[311] = exp_valid ? exp_out[311] : encrypted_data_buf[311];   // modexp_top.v(222)
    assign encrypted_data_buf_next[310] = exp_valid ? exp_out[310] : encrypted_data_buf[310];   // modexp_top.v(222)
    assign encrypted_data_buf_next[309] = exp_valid ? exp_out[309] : encrypted_data_buf[309];   // modexp_top.v(222)
    assign encrypted_data_buf_next[308] = exp_valid ? exp_out[308] : encrypted_data_buf[308];   // modexp_top.v(222)
    assign encrypted_data_buf_next[307] = exp_valid ? exp_out[307] : encrypted_data_buf[307];   // modexp_top.v(222)
    assign encrypted_data_buf_next[306] = exp_valid ? exp_out[306] : encrypted_data_buf[306];   // modexp_top.v(222)
    assign encrypted_data_buf_next[305] = exp_valid ? exp_out[305] : encrypted_data_buf[305];   // modexp_top.v(222)
    assign encrypted_data_buf_next[304] = exp_valid ? exp_out[304] : encrypted_data_buf[304];   // modexp_top.v(222)
    assign encrypted_data_buf_next[303] = exp_valid ? exp_out[303] : encrypted_data_buf[303];   // modexp_top.v(222)
    assign encrypted_data_buf_next[302] = exp_valid ? exp_out[302] : encrypted_data_buf[302];   // modexp_top.v(222)
    assign encrypted_data_buf_next[301] = exp_valid ? exp_out[301] : encrypted_data_buf[301];   // modexp_top.v(222)
    assign encrypted_data_buf_next[300] = exp_valid ? exp_out[300] : encrypted_data_buf[300];   // modexp_top.v(222)
    assign encrypted_data_buf_next[299] = exp_valid ? exp_out[299] : encrypted_data_buf[299];   // modexp_top.v(222)
    assign encrypted_data_buf_next[298] = exp_valid ? exp_out[298] : encrypted_data_buf[298];   // modexp_top.v(222)
    assign encrypted_data_buf_next[297] = exp_valid ? exp_out[297] : encrypted_data_buf[297];   // modexp_top.v(222)
    assign encrypted_data_buf_next[296] = exp_valid ? exp_out[296] : encrypted_data_buf[296];   // modexp_top.v(222)
    assign encrypted_data_buf_next[295] = exp_valid ? exp_out[295] : encrypted_data_buf[295];   // modexp_top.v(222)
    assign encrypted_data_buf_next[294] = exp_valid ? exp_out[294] : encrypted_data_buf[294];   // modexp_top.v(222)
    assign encrypted_data_buf_next[293] = exp_valid ? exp_out[293] : encrypted_data_buf[293];   // modexp_top.v(222)
    assign encrypted_data_buf_next[292] = exp_valid ? exp_out[292] : encrypted_data_buf[292];   // modexp_top.v(222)
    assign encrypted_data_buf_next[291] = exp_valid ? exp_out[291] : encrypted_data_buf[291];   // modexp_top.v(222)
    assign encrypted_data_buf_next[290] = exp_valid ? exp_out[290] : encrypted_data_buf[290];   // modexp_top.v(222)
    assign encrypted_data_buf_next[289] = exp_valid ? exp_out[289] : encrypted_data_buf[289];   // modexp_top.v(222)
    assign encrypted_data_buf_next[288] = exp_valid ? exp_out[288] : encrypted_data_buf[288];   // modexp_top.v(222)
    assign encrypted_data_buf_next[287] = exp_valid ? exp_out[287] : encrypted_data_buf[287];   // modexp_top.v(222)
    assign encrypted_data_buf_next[286] = exp_valid ? exp_out[286] : encrypted_data_buf[286];   // modexp_top.v(222)
    assign encrypted_data_buf_next[285] = exp_valid ? exp_out[285] : encrypted_data_buf[285];   // modexp_top.v(222)
    assign encrypted_data_buf_next[284] = exp_valid ? exp_out[284] : encrypted_data_buf[284];   // modexp_top.v(222)
    assign encrypted_data_buf_next[283] = exp_valid ? exp_out[283] : encrypted_data_buf[283];   // modexp_top.v(222)
    assign encrypted_data_buf_next[282] = exp_valid ? exp_out[282] : encrypted_data_buf[282];   // modexp_top.v(222)
    assign encrypted_data_buf_next[281] = exp_valid ? exp_out[281] : encrypted_data_buf[281];   // modexp_top.v(222)
    assign encrypted_data_buf_next[280] = exp_valid ? exp_out[280] : encrypted_data_buf[280];   // modexp_top.v(222)
    assign encrypted_data_buf_next[279] = exp_valid ? exp_out[279] : encrypted_data_buf[279];   // modexp_top.v(222)
    assign encrypted_data_buf_next[278] = exp_valid ? exp_out[278] : encrypted_data_buf[278];   // modexp_top.v(222)
    assign encrypted_data_buf_next[277] = exp_valid ? exp_out[277] : encrypted_data_buf[277];   // modexp_top.v(222)
    assign encrypted_data_buf_next[276] = exp_valid ? exp_out[276] : encrypted_data_buf[276];   // modexp_top.v(222)
    assign encrypted_data_buf_next[275] = exp_valid ? exp_out[275] : encrypted_data_buf[275];   // modexp_top.v(222)
    assign encrypted_data_buf_next[274] = exp_valid ? exp_out[274] : encrypted_data_buf[274];   // modexp_top.v(222)
    assign encrypted_data_buf_next[273] = exp_valid ? exp_out[273] : encrypted_data_buf[273];   // modexp_top.v(222)
    assign encrypted_data_buf_next[272] = exp_valid ? exp_out[272] : encrypted_data_buf[272];   // modexp_top.v(222)
    assign encrypted_data_buf_next[271] = exp_valid ? exp_out[271] : encrypted_data_buf[271];   // modexp_top.v(222)
    assign encrypted_data_buf_next[270] = exp_valid ? exp_out[270] : encrypted_data_buf[270];   // modexp_top.v(222)
    assign encrypted_data_buf_next[269] = exp_valid ? exp_out[269] : encrypted_data_buf[269];   // modexp_top.v(222)
    assign encrypted_data_buf_next[268] = exp_valid ? exp_out[268] : encrypted_data_buf[268];   // modexp_top.v(222)
    assign encrypted_data_buf_next[267] = exp_valid ? exp_out[267] : encrypted_data_buf[267];   // modexp_top.v(222)
    assign encrypted_data_buf_next[266] = exp_valid ? exp_out[266] : encrypted_data_buf[266];   // modexp_top.v(222)
    assign encrypted_data_buf_next[265] = exp_valid ? exp_out[265] : encrypted_data_buf[265];   // modexp_top.v(222)
    assign encrypted_data_buf_next[264] = exp_valid ? exp_out[264] : encrypted_data_buf[264];   // modexp_top.v(222)
    assign encrypted_data_buf_next[263] = exp_valid ? exp_out[263] : encrypted_data_buf[263];   // modexp_top.v(222)
    assign encrypted_data_buf_next[262] = exp_valid ? exp_out[262] : encrypted_data_buf[262];   // modexp_top.v(222)
    assign encrypted_data_buf_next[261] = exp_valid ? exp_out[261] : encrypted_data_buf[261];   // modexp_top.v(222)
    assign encrypted_data_buf_next[260] = exp_valid ? exp_out[260] : encrypted_data_buf[260];   // modexp_top.v(222)
    assign encrypted_data_buf_next[259] = exp_valid ? exp_out[259] : encrypted_data_buf[259];   // modexp_top.v(222)
    assign encrypted_data_buf_next[258] = exp_valid ? exp_out[258] : encrypted_data_buf[258];   // modexp_top.v(222)
    assign encrypted_data_buf_next[257] = exp_valid ? exp_out[257] : encrypted_data_buf[257];   // modexp_top.v(222)
    assign encrypted_data_buf_next[256] = exp_valid ? exp_out[256] : encrypted_data_buf[256];   // modexp_top.v(222)
    assign encrypted_data_buf_next[255] = exp_valid ? exp_out[255] : encrypted_data_buf[255];   // modexp_top.v(222)
    assign encrypted_data_buf_next[254] = exp_valid ? exp_out[254] : encrypted_data_buf[254];   // modexp_top.v(222)
    assign encrypted_data_buf_next[253] = exp_valid ? exp_out[253] : encrypted_data_buf[253];   // modexp_top.v(222)
    assign encrypted_data_buf_next[252] = exp_valid ? exp_out[252] : encrypted_data_buf[252];   // modexp_top.v(222)
    assign encrypted_data_buf_next[251] = exp_valid ? exp_out[251] : encrypted_data_buf[251];   // modexp_top.v(222)
    assign encrypted_data_buf_next[250] = exp_valid ? exp_out[250] : encrypted_data_buf[250];   // modexp_top.v(222)
    assign encrypted_data_buf_next[249] = exp_valid ? exp_out[249] : encrypted_data_buf[249];   // modexp_top.v(222)
    assign encrypted_data_buf_next[248] = exp_valid ? exp_out[248] : encrypted_data_buf[248];   // modexp_top.v(222)
    assign encrypted_data_buf_next[247] = exp_valid ? exp_out[247] : encrypted_data_buf[247];   // modexp_top.v(222)
    assign encrypted_data_buf_next[246] = exp_valid ? exp_out[246] : encrypted_data_buf[246];   // modexp_top.v(222)
    assign encrypted_data_buf_next[245] = exp_valid ? exp_out[245] : encrypted_data_buf[245];   // modexp_top.v(222)
    assign encrypted_data_buf_next[244] = exp_valid ? exp_out[244] : encrypted_data_buf[244];   // modexp_top.v(222)
    assign encrypted_data_buf_next[243] = exp_valid ? exp_out[243] : encrypted_data_buf[243];   // modexp_top.v(222)
    assign encrypted_data_buf_next[242] = exp_valid ? exp_out[242] : encrypted_data_buf[242];   // modexp_top.v(222)
    assign encrypted_data_buf_next[241] = exp_valid ? exp_out[241] : encrypted_data_buf[241];   // modexp_top.v(222)
    assign encrypted_data_buf_next[240] = exp_valid ? exp_out[240] : encrypted_data_buf[240];   // modexp_top.v(222)
    assign encrypted_data_buf_next[239] = exp_valid ? exp_out[239] : encrypted_data_buf[239];   // modexp_top.v(222)
    assign encrypted_data_buf_next[238] = exp_valid ? exp_out[238] : encrypted_data_buf[238];   // modexp_top.v(222)
    assign encrypted_data_buf_next[237] = exp_valid ? exp_out[237] : encrypted_data_buf[237];   // modexp_top.v(222)
    assign encrypted_data_buf_next[236] = exp_valid ? exp_out[236] : encrypted_data_buf[236];   // modexp_top.v(222)
    assign encrypted_data_buf_next[235] = exp_valid ? exp_out[235] : encrypted_data_buf[235];   // modexp_top.v(222)
    assign encrypted_data_buf_next[234] = exp_valid ? exp_out[234] : encrypted_data_buf[234];   // modexp_top.v(222)
    assign encrypted_data_buf_next[233] = exp_valid ? exp_out[233] : encrypted_data_buf[233];   // modexp_top.v(222)
    assign encrypted_data_buf_next[232] = exp_valid ? exp_out[232] : encrypted_data_buf[232];   // modexp_top.v(222)
    assign encrypted_data_buf_next[231] = exp_valid ? exp_out[231] : encrypted_data_buf[231];   // modexp_top.v(222)
    assign encrypted_data_buf_next[230] = exp_valid ? exp_out[230] : encrypted_data_buf[230];   // modexp_top.v(222)
    assign encrypted_data_buf_next[229] = exp_valid ? exp_out[229] : encrypted_data_buf[229];   // modexp_top.v(222)
    assign encrypted_data_buf_next[228] = exp_valid ? exp_out[228] : encrypted_data_buf[228];   // modexp_top.v(222)
    assign encrypted_data_buf_next[227] = exp_valid ? exp_out[227] : encrypted_data_buf[227];   // modexp_top.v(222)
    assign encrypted_data_buf_next[226] = exp_valid ? exp_out[226] : encrypted_data_buf[226];   // modexp_top.v(222)
    assign encrypted_data_buf_next[225] = exp_valid ? exp_out[225] : encrypted_data_buf[225];   // modexp_top.v(222)
    assign encrypted_data_buf_next[224] = exp_valid ? exp_out[224] : encrypted_data_buf[224];   // modexp_top.v(222)
    assign encrypted_data_buf_next[223] = exp_valid ? exp_out[223] : encrypted_data_buf[223];   // modexp_top.v(222)
    assign encrypted_data_buf_next[222] = exp_valid ? exp_out[222] : encrypted_data_buf[222];   // modexp_top.v(222)
    assign encrypted_data_buf_next[221] = exp_valid ? exp_out[221] : encrypted_data_buf[221];   // modexp_top.v(222)
    assign encrypted_data_buf_next[220] = exp_valid ? exp_out[220] : encrypted_data_buf[220];   // modexp_top.v(222)
    assign encrypted_data_buf_next[219] = exp_valid ? exp_out[219] : encrypted_data_buf[219];   // modexp_top.v(222)
    assign encrypted_data_buf_next[218] = exp_valid ? exp_out[218] : encrypted_data_buf[218];   // modexp_top.v(222)
    assign encrypted_data_buf_next[217] = exp_valid ? exp_out[217] : encrypted_data_buf[217];   // modexp_top.v(222)
    assign encrypted_data_buf_next[216] = exp_valid ? exp_out[216] : encrypted_data_buf[216];   // modexp_top.v(222)
    assign encrypted_data_buf_next[215] = exp_valid ? exp_out[215] : encrypted_data_buf[215];   // modexp_top.v(222)
    assign encrypted_data_buf_next[214] = exp_valid ? exp_out[214] : encrypted_data_buf[214];   // modexp_top.v(222)
    assign encrypted_data_buf_next[213] = exp_valid ? exp_out[213] : encrypted_data_buf[213];   // modexp_top.v(222)
    assign encrypted_data_buf_next[212] = exp_valid ? exp_out[212] : encrypted_data_buf[212];   // modexp_top.v(222)
    assign encrypted_data_buf_next[211] = exp_valid ? exp_out[211] : encrypted_data_buf[211];   // modexp_top.v(222)
    assign encrypted_data_buf_next[210] = exp_valid ? exp_out[210] : encrypted_data_buf[210];   // modexp_top.v(222)
    assign encrypted_data_buf_next[209] = exp_valid ? exp_out[209] : encrypted_data_buf[209];   // modexp_top.v(222)
    assign encrypted_data_buf_next[208] = exp_valid ? exp_out[208] : encrypted_data_buf[208];   // modexp_top.v(222)
    assign encrypted_data_buf_next[207] = exp_valid ? exp_out[207] : encrypted_data_buf[207];   // modexp_top.v(222)
    assign encrypted_data_buf_next[206] = exp_valid ? exp_out[206] : encrypted_data_buf[206];   // modexp_top.v(222)
    assign encrypted_data_buf_next[205] = exp_valid ? exp_out[205] : encrypted_data_buf[205];   // modexp_top.v(222)
    assign encrypted_data_buf_next[204] = exp_valid ? exp_out[204] : encrypted_data_buf[204];   // modexp_top.v(222)
    assign encrypted_data_buf_next[203] = exp_valid ? exp_out[203] : encrypted_data_buf[203];   // modexp_top.v(222)
    assign encrypted_data_buf_next[202] = exp_valid ? exp_out[202] : encrypted_data_buf[202];   // modexp_top.v(222)
    assign encrypted_data_buf_next[201] = exp_valid ? exp_out[201] : encrypted_data_buf[201];   // modexp_top.v(222)
    assign encrypted_data_buf_next[200] = exp_valid ? exp_out[200] : encrypted_data_buf[200];   // modexp_top.v(222)
    assign encrypted_data_buf_next[199] = exp_valid ? exp_out[199] : encrypted_data_buf[199];   // modexp_top.v(222)
    assign encrypted_data_buf_next[198] = exp_valid ? exp_out[198] : encrypted_data_buf[198];   // modexp_top.v(222)
    assign encrypted_data_buf_next[197] = exp_valid ? exp_out[197] : encrypted_data_buf[197];   // modexp_top.v(222)
    assign encrypted_data_buf_next[196] = exp_valid ? exp_out[196] : encrypted_data_buf[196];   // modexp_top.v(222)
    assign encrypted_data_buf_next[195] = exp_valid ? exp_out[195] : encrypted_data_buf[195];   // modexp_top.v(222)
    assign encrypted_data_buf_next[194] = exp_valid ? exp_out[194] : encrypted_data_buf[194];   // modexp_top.v(222)
    assign encrypted_data_buf_next[193] = exp_valid ? exp_out[193] : encrypted_data_buf[193];   // modexp_top.v(222)
    assign encrypted_data_buf_next[192] = exp_valid ? exp_out[192] : encrypted_data_buf[192];   // modexp_top.v(222)
    assign encrypted_data_buf_next[191] = exp_valid ? exp_out[191] : encrypted_data_buf[191];   // modexp_top.v(222)
    assign encrypted_data_buf_next[190] = exp_valid ? exp_out[190] : encrypted_data_buf[190];   // modexp_top.v(222)
    assign encrypted_data_buf_next[189] = exp_valid ? exp_out[189] : encrypted_data_buf[189];   // modexp_top.v(222)
    assign encrypted_data_buf_next[188] = exp_valid ? exp_out[188] : encrypted_data_buf[188];   // modexp_top.v(222)
    assign encrypted_data_buf_next[187] = exp_valid ? exp_out[187] : encrypted_data_buf[187];   // modexp_top.v(222)
    assign encrypted_data_buf_next[186] = exp_valid ? exp_out[186] : encrypted_data_buf[186];   // modexp_top.v(222)
    assign encrypted_data_buf_next[185] = exp_valid ? exp_out[185] : encrypted_data_buf[185];   // modexp_top.v(222)
    assign encrypted_data_buf_next[184] = exp_valid ? exp_out[184] : encrypted_data_buf[184];   // modexp_top.v(222)
    assign encrypted_data_buf_next[183] = exp_valid ? exp_out[183] : encrypted_data_buf[183];   // modexp_top.v(222)
    assign encrypted_data_buf_next[182] = exp_valid ? exp_out[182] : encrypted_data_buf[182];   // modexp_top.v(222)
    assign encrypted_data_buf_next[181] = exp_valid ? exp_out[181] : encrypted_data_buf[181];   // modexp_top.v(222)
    assign encrypted_data_buf_next[180] = exp_valid ? exp_out[180] : encrypted_data_buf[180];   // modexp_top.v(222)
    assign encrypted_data_buf_next[179] = exp_valid ? exp_out[179] : encrypted_data_buf[179];   // modexp_top.v(222)
    assign encrypted_data_buf_next[178] = exp_valid ? exp_out[178] : encrypted_data_buf[178];   // modexp_top.v(222)
    assign encrypted_data_buf_next[177] = exp_valid ? exp_out[177] : encrypted_data_buf[177];   // modexp_top.v(222)
    assign encrypted_data_buf_next[176] = exp_valid ? exp_out[176] : encrypted_data_buf[176];   // modexp_top.v(222)
    assign encrypted_data_buf_next[175] = exp_valid ? exp_out[175] : encrypted_data_buf[175];   // modexp_top.v(222)
    assign encrypted_data_buf_next[174] = exp_valid ? exp_out[174] : encrypted_data_buf[174];   // modexp_top.v(222)
    assign encrypted_data_buf_next[173] = exp_valid ? exp_out[173] : encrypted_data_buf[173];   // modexp_top.v(222)
    assign encrypted_data_buf_next[172] = exp_valid ? exp_out[172] : encrypted_data_buf[172];   // modexp_top.v(222)
    assign encrypted_data_buf_next[171] = exp_valid ? exp_out[171] : encrypted_data_buf[171];   // modexp_top.v(222)
    assign encrypted_data_buf_next[170] = exp_valid ? exp_out[170] : encrypted_data_buf[170];   // modexp_top.v(222)
    assign encrypted_data_buf_next[169] = exp_valid ? exp_out[169] : encrypted_data_buf[169];   // modexp_top.v(222)
    assign encrypted_data_buf_next[168] = exp_valid ? exp_out[168] : encrypted_data_buf[168];   // modexp_top.v(222)
    assign encrypted_data_buf_next[167] = exp_valid ? exp_out[167] : encrypted_data_buf[167];   // modexp_top.v(222)
    assign encrypted_data_buf_next[166] = exp_valid ? exp_out[166] : encrypted_data_buf[166];   // modexp_top.v(222)
    assign encrypted_data_buf_next[165] = exp_valid ? exp_out[165] : encrypted_data_buf[165];   // modexp_top.v(222)
    assign encrypted_data_buf_next[164] = exp_valid ? exp_out[164] : encrypted_data_buf[164];   // modexp_top.v(222)
    assign encrypted_data_buf_next[163] = exp_valid ? exp_out[163] : encrypted_data_buf[163];   // modexp_top.v(222)
    assign encrypted_data_buf_next[162] = exp_valid ? exp_out[162] : encrypted_data_buf[162];   // modexp_top.v(222)
    assign encrypted_data_buf_next[161] = exp_valid ? exp_out[161] : encrypted_data_buf[161];   // modexp_top.v(222)
    assign encrypted_data_buf_next[160] = exp_valid ? exp_out[160] : encrypted_data_buf[160];   // modexp_top.v(222)
    assign encrypted_data_buf_next[159] = exp_valid ? exp_out[159] : encrypted_data_buf[159];   // modexp_top.v(222)
    assign encrypted_data_buf_next[158] = exp_valid ? exp_out[158] : encrypted_data_buf[158];   // modexp_top.v(222)
    assign encrypted_data_buf_next[157] = exp_valid ? exp_out[157] : encrypted_data_buf[157];   // modexp_top.v(222)
    assign encrypted_data_buf_next[156] = exp_valid ? exp_out[156] : encrypted_data_buf[156];   // modexp_top.v(222)
    assign encrypted_data_buf_next[155] = exp_valid ? exp_out[155] : encrypted_data_buf[155];   // modexp_top.v(222)
    assign encrypted_data_buf_next[154] = exp_valid ? exp_out[154] : encrypted_data_buf[154];   // modexp_top.v(222)
    assign encrypted_data_buf_next[153] = exp_valid ? exp_out[153] : encrypted_data_buf[153];   // modexp_top.v(222)
    assign encrypted_data_buf_next[152] = exp_valid ? exp_out[152] : encrypted_data_buf[152];   // modexp_top.v(222)
    assign encrypted_data_buf_next[151] = exp_valid ? exp_out[151] : encrypted_data_buf[151];   // modexp_top.v(222)
    assign encrypted_data_buf_next[150] = exp_valid ? exp_out[150] : encrypted_data_buf[150];   // modexp_top.v(222)
    assign encrypted_data_buf_next[149] = exp_valid ? exp_out[149] : encrypted_data_buf[149];   // modexp_top.v(222)
    assign encrypted_data_buf_next[148] = exp_valid ? exp_out[148] : encrypted_data_buf[148];   // modexp_top.v(222)
    assign encrypted_data_buf_next[147] = exp_valid ? exp_out[147] : encrypted_data_buf[147];   // modexp_top.v(222)
    assign encrypted_data_buf_next[146] = exp_valid ? exp_out[146] : encrypted_data_buf[146];   // modexp_top.v(222)
    assign encrypted_data_buf_next[145] = exp_valid ? exp_out[145] : encrypted_data_buf[145];   // modexp_top.v(222)
    assign encrypted_data_buf_next[144] = exp_valid ? exp_out[144] : encrypted_data_buf[144];   // modexp_top.v(222)
    assign encrypted_data_buf_next[143] = exp_valid ? exp_out[143] : encrypted_data_buf[143];   // modexp_top.v(222)
    assign encrypted_data_buf_next[142] = exp_valid ? exp_out[142] : encrypted_data_buf[142];   // modexp_top.v(222)
    assign encrypted_data_buf_next[141] = exp_valid ? exp_out[141] : encrypted_data_buf[141];   // modexp_top.v(222)
    assign encrypted_data_buf_next[140] = exp_valid ? exp_out[140] : encrypted_data_buf[140];   // modexp_top.v(222)
    assign encrypted_data_buf_next[139] = exp_valid ? exp_out[139] : encrypted_data_buf[139];   // modexp_top.v(222)
    assign encrypted_data_buf_next[138] = exp_valid ? exp_out[138] : encrypted_data_buf[138];   // modexp_top.v(222)
    assign encrypted_data_buf_next[137] = exp_valid ? exp_out[137] : encrypted_data_buf[137];   // modexp_top.v(222)
    assign encrypted_data_buf_next[136] = exp_valid ? exp_out[136] : encrypted_data_buf[136];   // modexp_top.v(222)
    assign encrypted_data_buf_next[135] = exp_valid ? exp_out[135] : encrypted_data_buf[135];   // modexp_top.v(222)
    assign encrypted_data_buf_next[134] = exp_valid ? exp_out[134] : encrypted_data_buf[134];   // modexp_top.v(222)
    assign encrypted_data_buf_next[133] = exp_valid ? exp_out[133] : encrypted_data_buf[133];   // modexp_top.v(222)
    assign encrypted_data_buf_next[132] = exp_valid ? exp_out[132] : encrypted_data_buf[132];   // modexp_top.v(222)
    assign encrypted_data_buf_next[131] = exp_valid ? exp_out[131] : encrypted_data_buf[131];   // modexp_top.v(222)
    assign encrypted_data_buf_next[130] = exp_valid ? exp_out[130] : encrypted_data_buf[130];   // modexp_top.v(222)
    assign encrypted_data_buf_next[129] = exp_valid ? exp_out[129] : encrypted_data_buf[129];   // modexp_top.v(222)
    assign encrypted_data_buf_next[128] = exp_valid ? exp_out[128] : encrypted_data_buf[128];   // modexp_top.v(222)
    assign encrypted_data_buf_next[127] = exp_valid ? exp_out[127] : encrypted_data_buf[127];   // modexp_top.v(222)
    assign encrypted_data_buf_next[126] = exp_valid ? exp_out[126] : encrypted_data_buf[126];   // modexp_top.v(222)
    assign encrypted_data_buf_next[125] = exp_valid ? exp_out[125] : encrypted_data_buf[125];   // modexp_top.v(222)
    assign encrypted_data_buf_next[124] = exp_valid ? exp_out[124] : encrypted_data_buf[124];   // modexp_top.v(222)
    assign encrypted_data_buf_next[123] = exp_valid ? exp_out[123] : encrypted_data_buf[123];   // modexp_top.v(222)
    assign encrypted_data_buf_next[122] = exp_valid ? exp_out[122] : encrypted_data_buf[122];   // modexp_top.v(222)
    assign encrypted_data_buf_next[121] = exp_valid ? exp_out[121] : encrypted_data_buf[121];   // modexp_top.v(222)
    assign encrypted_data_buf_next[120] = exp_valid ? exp_out[120] : encrypted_data_buf[120];   // modexp_top.v(222)
    assign encrypted_data_buf_next[119] = exp_valid ? exp_out[119] : encrypted_data_buf[119];   // modexp_top.v(222)
    assign encrypted_data_buf_next[118] = exp_valid ? exp_out[118] : encrypted_data_buf[118];   // modexp_top.v(222)
    assign encrypted_data_buf_next[117] = exp_valid ? exp_out[117] : encrypted_data_buf[117];   // modexp_top.v(222)
    assign encrypted_data_buf_next[116] = exp_valid ? exp_out[116] : encrypted_data_buf[116];   // modexp_top.v(222)
    assign encrypted_data_buf_next[115] = exp_valid ? exp_out[115] : encrypted_data_buf[115];   // modexp_top.v(222)
    assign encrypted_data_buf_next[114] = exp_valid ? exp_out[114] : encrypted_data_buf[114];   // modexp_top.v(222)
    assign encrypted_data_buf_next[113] = exp_valid ? exp_out[113] : encrypted_data_buf[113];   // modexp_top.v(222)
    assign encrypted_data_buf_next[112] = exp_valid ? exp_out[112] : encrypted_data_buf[112];   // modexp_top.v(222)
    assign encrypted_data_buf_next[111] = exp_valid ? exp_out[111] : encrypted_data_buf[111];   // modexp_top.v(222)
    assign encrypted_data_buf_next[110] = exp_valid ? exp_out[110] : encrypted_data_buf[110];   // modexp_top.v(222)
    assign encrypted_data_buf_next[109] = exp_valid ? exp_out[109] : encrypted_data_buf[109];   // modexp_top.v(222)
    assign encrypted_data_buf_next[108] = exp_valid ? exp_out[108] : encrypted_data_buf[108];   // modexp_top.v(222)
    assign encrypted_data_buf_next[107] = exp_valid ? exp_out[107] : encrypted_data_buf[107];   // modexp_top.v(222)
    assign encrypted_data_buf_next[106] = exp_valid ? exp_out[106] : encrypted_data_buf[106];   // modexp_top.v(222)
    assign encrypted_data_buf_next[105] = exp_valid ? exp_out[105] : encrypted_data_buf[105];   // modexp_top.v(222)
    assign encrypted_data_buf_next[104] = exp_valid ? exp_out[104] : encrypted_data_buf[104];   // modexp_top.v(222)
    assign encrypted_data_buf_next[103] = exp_valid ? exp_out[103] : encrypted_data_buf[103];   // modexp_top.v(222)
    assign encrypted_data_buf_next[102] = exp_valid ? exp_out[102] : encrypted_data_buf[102];   // modexp_top.v(222)
    assign encrypted_data_buf_next[101] = exp_valid ? exp_out[101] : encrypted_data_buf[101];   // modexp_top.v(222)
    assign encrypted_data_buf_next[100] = exp_valid ? exp_out[100] : encrypted_data_buf[100];   // modexp_top.v(222)
    assign encrypted_data_buf_next[99] = exp_valid ? exp_out[99] : encrypted_data_buf[99];   // modexp_top.v(222)
    assign encrypted_data_buf_next[98] = exp_valid ? exp_out[98] : encrypted_data_buf[98];   // modexp_top.v(222)
    assign encrypted_data_buf_next[97] = exp_valid ? exp_out[97] : encrypted_data_buf[97];   // modexp_top.v(222)
    assign encrypted_data_buf_next[96] = exp_valid ? exp_out[96] : encrypted_data_buf[96];   // modexp_top.v(222)
    assign encrypted_data_buf_next[95] = exp_valid ? exp_out[95] : encrypted_data_buf[95];   // modexp_top.v(222)
    assign encrypted_data_buf_next[94] = exp_valid ? exp_out[94] : encrypted_data_buf[94];   // modexp_top.v(222)
    assign encrypted_data_buf_next[93] = exp_valid ? exp_out[93] : encrypted_data_buf[93];   // modexp_top.v(222)
    assign encrypted_data_buf_next[92] = exp_valid ? exp_out[92] : encrypted_data_buf[92];   // modexp_top.v(222)
    assign encrypted_data_buf_next[91] = exp_valid ? exp_out[91] : encrypted_data_buf[91];   // modexp_top.v(222)
    assign encrypted_data_buf_next[90] = exp_valid ? exp_out[90] : encrypted_data_buf[90];   // modexp_top.v(222)
    assign encrypted_data_buf_next[89] = exp_valid ? exp_out[89] : encrypted_data_buf[89];   // modexp_top.v(222)
    assign encrypted_data_buf_next[88] = exp_valid ? exp_out[88] : encrypted_data_buf[88];   // modexp_top.v(222)
    assign encrypted_data_buf_next[87] = exp_valid ? exp_out[87] : encrypted_data_buf[87];   // modexp_top.v(222)
    assign encrypted_data_buf_next[86] = exp_valid ? exp_out[86] : encrypted_data_buf[86];   // modexp_top.v(222)
    assign encrypted_data_buf_next[85] = exp_valid ? exp_out[85] : encrypted_data_buf[85];   // modexp_top.v(222)
    assign encrypted_data_buf_next[84] = exp_valid ? exp_out[84] : encrypted_data_buf[84];   // modexp_top.v(222)
    assign encrypted_data_buf_next[83] = exp_valid ? exp_out[83] : encrypted_data_buf[83];   // modexp_top.v(222)
    assign encrypted_data_buf_next[82] = exp_valid ? exp_out[82] : encrypted_data_buf[82];   // modexp_top.v(222)
    assign encrypted_data_buf_next[81] = exp_valid ? exp_out[81] : encrypted_data_buf[81];   // modexp_top.v(222)
    assign encrypted_data_buf_next[80] = exp_valid ? exp_out[80] : encrypted_data_buf[80];   // modexp_top.v(222)
    assign encrypted_data_buf_next[79] = exp_valid ? exp_out[79] : encrypted_data_buf[79];   // modexp_top.v(222)
    assign encrypted_data_buf_next[78] = exp_valid ? exp_out[78] : encrypted_data_buf[78];   // modexp_top.v(222)
    assign encrypted_data_buf_next[77] = exp_valid ? exp_out[77] : encrypted_data_buf[77];   // modexp_top.v(222)
    assign encrypted_data_buf_next[76] = exp_valid ? exp_out[76] : encrypted_data_buf[76];   // modexp_top.v(222)
    assign encrypted_data_buf_next[75] = exp_valid ? exp_out[75] : encrypted_data_buf[75];   // modexp_top.v(222)
    assign encrypted_data_buf_next[74] = exp_valid ? exp_out[74] : encrypted_data_buf[74];   // modexp_top.v(222)
    assign encrypted_data_buf_next[73] = exp_valid ? exp_out[73] : encrypted_data_buf[73];   // modexp_top.v(222)
    assign encrypted_data_buf_next[72] = exp_valid ? exp_out[72] : encrypted_data_buf[72];   // modexp_top.v(222)
    assign encrypted_data_buf_next[71] = exp_valid ? exp_out[71] : encrypted_data_buf[71];   // modexp_top.v(222)
    assign encrypted_data_buf_next[70] = exp_valid ? exp_out[70] : encrypted_data_buf[70];   // modexp_top.v(222)
    assign encrypted_data_buf_next[69] = exp_valid ? exp_out[69] : encrypted_data_buf[69];   // modexp_top.v(222)
    assign encrypted_data_buf_next[68] = exp_valid ? exp_out[68] : encrypted_data_buf[68];   // modexp_top.v(222)
    assign encrypted_data_buf_next[67] = exp_valid ? exp_out[67] : encrypted_data_buf[67];   // modexp_top.v(222)
    assign encrypted_data_buf_next[66] = exp_valid ? exp_out[66] : encrypted_data_buf[66];   // modexp_top.v(222)
    assign encrypted_data_buf_next[65] = exp_valid ? exp_out[65] : encrypted_data_buf[65];   // modexp_top.v(222)
    assign encrypted_data_buf_next[64] = exp_valid ? exp_out[64] : encrypted_data_buf[64];   // modexp_top.v(222)
    assign encrypted_data_buf_next[63] = exp_valid ? exp_out[63] : encrypted_data_buf[63];   // modexp_top.v(222)
    assign encrypted_data_buf_next[62] = exp_valid ? exp_out[62] : encrypted_data_buf[62];   // modexp_top.v(222)
    assign encrypted_data_buf_next[61] = exp_valid ? exp_out[61] : encrypted_data_buf[61];   // modexp_top.v(222)
    assign encrypted_data_buf_next[60] = exp_valid ? exp_out[60] : encrypted_data_buf[60];   // modexp_top.v(222)
    assign encrypted_data_buf_next[59] = exp_valid ? exp_out[59] : encrypted_data_buf[59];   // modexp_top.v(222)
    assign encrypted_data_buf_next[58] = exp_valid ? exp_out[58] : encrypted_data_buf[58];   // modexp_top.v(222)
    assign encrypted_data_buf_next[57] = exp_valid ? exp_out[57] : encrypted_data_buf[57];   // modexp_top.v(222)
    assign encrypted_data_buf_next[56] = exp_valid ? exp_out[56] : encrypted_data_buf[56];   // modexp_top.v(222)
    assign encrypted_data_buf_next[55] = exp_valid ? exp_out[55] : encrypted_data_buf[55];   // modexp_top.v(222)
    assign encrypted_data_buf_next[54] = exp_valid ? exp_out[54] : encrypted_data_buf[54];   // modexp_top.v(222)
    assign encrypted_data_buf_next[53] = exp_valid ? exp_out[53] : encrypted_data_buf[53];   // modexp_top.v(222)
    assign encrypted_data_buf_next[52] = exp_valid ? exp_out[52] : encrypted_data_buf[52];   // modexp_top.v(222)
    assign encrypted_data_buf_next[51] = exp_valid ? exp_out[51] : encrypted_data_buf[51];   // modexp_top.v(222)
    assign encrypted_data_buf_next[50] = exp_valid ? exp_out[50] : encrypted_data_buf[50];   // modexp_top.v(222)
    assign encrypted_data_buf_next[49] = exp_valid ? exp_out[49] : encrypted_data_buf[49];   // modexp_top.v(222)
    assign encrypted_data_buf_next[48] = exp_valid ? exp_out[48] : encrypted_data_buf[48];   // modexp_top.v(222)
    assign encrypted_data_buf_next[47] = exp_valid ? exp_out[47] : encrypted_data_buf[47];   // modexp_top.v(222)
    assign encrypted_data_buf_next[46] = exp_valid ? exp_out[46] : encrypted_data_buf[46];   // modexp_top.v(222)
    assign encrypted_data_buf_next[45] = exp_valid ? exp_out[45] : encrypted_data_buf[45];   // modexp_top.v(222)
    assign encrypted_data_buf_next[44] = exp_valid ? exp_out[44] : encrypted_data_buf[44];   // modexp_top.v(222)
    assign encrypted_data_buf_next[43] = exp_valid ? exp_out[43] : encrypted_data_buf[43];   // modexp_top.v(222)
    assign encrypted_data_buf_next[42] = exp_valid ? exp_out[42] : encrypted_data_buf[42];   // modexp_top.v(222)
    assign encrypted_data_buf_next[41] = exp_valid ? exp_out[41] : encrypted_data_buf[41];   // modexp_top.v(222)
    assign encrypted_data_buf_next[40] = exp_valid ? exp_out[40] : encrypted_data_buf[40];   // modexp_top.v(222)
    assign encrypted_data_buf_next[39] = exp_valid ? exp_out[39] : encrypted_data_buf[39];   // modexp_top.v(222)
    assign encrypted_data_buf_next[38] = exp_valid ? exp_out[38] : encrypted_data_buf[38];   // modexp_top.v(222)
    assign encrypted_data_buf_next[37] = exp_valid ? exp_out[37] : encrypted_data_buf[37];   // modexp_top.v(222)
    assign encrypted_data_buf_next[36] = exp_valid ? exp_out[36] : encrypted_data_buf[36];   // modexp_top.v(222)
    assign encrypted_data_buf_next[35] = exp_valid ? exp_out[35] : encrypted_data_buf[35];   // modexp_top.v(222)
    assign encrypted_data_buf_next[34] = exp_valid ? exp_out[34] : encrypted_data_buf[34];   // modexp_top.v(222)
    assign encrypted_data_buf_next[33] = exp_valid ? exp_out[33] : encrypted_data_buf[33];   // modexp_top.v(222)
    assign encrypted_data_buf_next[32] = exp_valid ? exp_out[32] : encrypted_data_buf[32];   // modexp_top.v(222)
    assign encrypted_data_buf_next[31] = exp_valid ? exp_out[31] : encrypted_data_buf[31];   // modexp_top.v(222)
    assign encrypted_data_buf_next[30] = exp_valid ? exp_out[30] : encrypted_data_buf[30];   // modexp_top.v(222)
    assign encrypted_data_buf_next[29] = exp_valid ? exp_out[29] : encrypted_data_buf[29];   // modexp_top.v(222)
    assign encrypted_data_buf_next[28] = exp_valid ? exp_out[28] : encrypted_data_buf[28];   // modexp_top.v(222)
    assign encrypted_data_buf_next[27] = exp_valid ? exp_out[27] : encrypted_data_buf[27];   // modexp_top.v(222)
    assign encrypted_data_buf_next[26] = exp_valid ? exp_out[26] : encrypted_data_buf[26];   // modexp_top.v(222)
    assign encrypted_data_buf_next[25] = exp_valid ? exp_out[25] : encrypted_data_buf[25];   // modexp_top.v(222)
    assign encrypted_data_buf_next[24] = exp_valid ? exp_out[24] : encrypted_data_buf[24];   // modexp_top.v(222)
    assign encrypted_data_buf_next[23] = exp_valid ? exp_out[23] : encrypted_data_buf[23];   // modexp_top.v(222)
    assign encrypted_data_buf_next[22] = exp_valid ? exp_out[22] : encrypted_data_buf[22];   // modexp_top.v(222)
    assign encrypted_data_buf_next[21] = exp_valid ? exp_out[21] : encrypted_data_buf[21];   // modexp_top.v(222)
    assign encrypted_data_buf_next[20] = exp_valid ? exp_out[20] : encrypted_data_buf[20];   // modexp_top.v(222)
    assign encrypted_data_buf_next[19] = exp_valid ? exp_out[19] : encrypted_data_buf[19];   // modexp_top.v(222)
    assign encrypted_data_buf_next[18] = exp_valid ? exp_out[18] : encrypted_data_buf[18];   // modexp_top.v(222)
    assign encrypted_data_buf_next[17] = exp_valid ? exp_out[17] : encrypted_data_buf[17];   // modexp_top.v(222)
    assign encrypted_data_buf_next[16] = exp_valid ? exp_out[16] : encrypted_data_buf[16];   // modexp_top.v(222)
    assign encrypted_data_buf_next[15] = exp_valid ? exp_out[15] : encrypted_data_buf[15];   // modexp_top.v(222)
    assign encrypted_data_buf_next[14] = exp_valid ? exp_out[14] : encrypted_data_buf[14];   // modexp_top.v(222)
    assign encrypted_data_buf_next[13] = exp_valid ? exp_out[13] : encrypted_data_buf[13];   // modexp_top.v(222)
    assign encrypted_data_buf_next[12] = exp_valid ? exp_out[12] : encrypted_data_buf[12];   // modexp_top.v(222)
    assign encrypted_data_buf_next[11] = exp_valid ? exp_out[11] : encrypted_data_buf[11];   // modexp_top.v(222)
    assign encrypted_data_buf_next[10] = exp_valid ? exp_out[10] : encrypted_data_buf[10];   // modexp_top.v(222)
    assign encrypted_data_buf_next[9] = exp_valid ? exp_out[9] : encrypted_data_buf[9];   // modexp_top.v(222)
    assign encrypted_data_buf_next[8] = exp_valid ? exp_out[8] : encrypted_data_buf[8];   // modexp_top.v(222)
    assign encrypted_data_buf_next[7] = exp_valid ? exp_out[7] : encrypted_data_buf[7];   // modexp_top.v(222)
    assign encrypted_data_buf_next[6] = exp_valid ? exp_out[6] : encrypted_data_buf[6];   // modexp_top.v(222)
    assign encrypted_data_buf_next[5] = exp_valid ? exp_out[5] : encrypted_data_buf[5];   // modexp_top.v(222)
    assign encrypted_data_buf_next[4] = exp_valid ? exp_out[4] : encrypted_data_buf[4];   // modexp_top.v(222)
    assign encrypted_data_buf_next[3] = exp_valid ? exp_out[3] : encrypted_data_buf[3];   // modexp_top.v(222)
    assign encrypted_data_buf_next[2] = exp_valid ? exp_out[2] : encrypted_data_buf[2];   // modexp_top.v(222)
    assign encrypted_data_buf_next[1] = exp_valid ? exp_out[1] : encrypted_data_buf[1];   // modexp_top.v(222)
    assign encrypted_data_buf_next[0] = exp_valid ? exp_out[0] : encrypted_data_buf[0];   // modexp_top.v(222)
    nor (n2254, n153, n152, n151, n150, n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(227)
    nor (n2262, n153, n152, n151, n150, n149, n148, byte_counter[1], 
        n146) ;   // modexp_top.v(228)
    nor (n2269, n153, n152, n151, n150, n149, n148, byte_counter[1], 
        byte_counter[0]) ;   // modexp_top.v(229)
    nor (n2277, n153, n152, n151, n150, n149, byte_counter[2], 
        n147, n146) ;   // modexp_top.v(230)
    nor (n2284, n153, n152, n151, n150, n149, byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(231)
    nor (n2291, n153, n152, n151, n150, n149, byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(232)
    nor (n2297, n153, n152, n151, n150, n149, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(233)
    nor (n2305, n153, n152, n151, n150, byte_counter[3], n148, 
        n147, n146) ;   // modexp_top.v(234)
    nor (n2312, n153, n152, n151, n150, byte_counter[3], n148, 
        n147, byte_counter[0]) ;   // modexp_top.v(235)
    nor (n2319, n153, n152, n151, n150, byte_counter[3], n148, 
        byte_counter[1], n146) ;   // modexp_top.v(236)
    nor (n2325, n153, n152, n151, n150, byte_counter[3], n148, 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(237)
    nor (n2332, n153, n152, n151, n150, byte_counter[3], byte_counter[2], 
        n147, n146) ;   // modexp_top.v(238)
    nor (n2338, n153, n152, n151, n150, byte_counter[3], byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(239)
    nor (n2344, n153, n152, n151, n150, byte_counter[3], byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(240)
    nor (n2349, n153, n152, n151, n150, byte_counter[3], byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(241)
    nor (n2357, n153, n152, n151, byte_counter[4], n149, n148, 
        n147, n146) ;   // modexp_top.v(242)
    nor (n2364, n153, n152, n151, byte_counter[4], n149, n148, 
        n147, byte_counter[0]) ;   // modexp_top.v(243)
    nor (n2371, n153, n152, n151, byte_counter[4], n149, n148, 
        byte_counter[1], n146) ;   // modexp_top.v(244)
    nor (n2377, n153, n152, n151, byte_counter[4], n149, n148, 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(245)
    nor (n2384, n153, n152, n151, byte_counter[4], n149, byte_counter[2], 
        n147, n146) ;   // modexp_top.v(246)
    nor (n2390, n153, n152, n151, byte_counter[4], n149, byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(247)
    nor (n2396, n153, n152, n151, byte_counter[4], n149, byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(248)
    nor (n2401, n153, n152, n151, byte_counter[4], n149, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(249)
    nor (n2408, n153, n152, n151, byte_counter[4], byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(250)
    nor (n2414, n153, n152, n151, byte_counter[4], byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(251)
    nor (n2420, n153, n152, n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(252)
    nor (n2425, n153, n152, n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(253)
    nor (n2431, n153, n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(254)
    nor (n2436, n153, n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(255)
    nor (n2441, n153, n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(256)
    nor (n2445, n153, n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(257)
    nor (n2453, n153, n152, byte_counter[5], n150, n149, n148, 
        n147, n146) ;   // modexp_top.v(258)
    nor (n2460, n153, n152, byte_counter[5], n150, n149, n148, 
        n147, byte_counter[0]) ;   // modexp_top.v(259)
    nor (n2467, n153, n152, byte_counter[5], n150, n149, n148, 
        byte_counter[1], n146) ;   // modexp_top.v(260)
    nor (n2473, n153, n152, byte_counter[5], n150, n149, n148, 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(261)
    nor (n2480, n153, n152, byte_counter[5], n150, n149, byte_counter[2], 
        n147, n146) ;   // modexp_top.v(262)
    nor (n2486, n153, n152, byte_counter[5], n150, n149, byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(263)
    nor (n2492, n153, n152, byte_counter[5], n150, n149, byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(264)
    nor (n2497, n153, n152, byte_counter[5], n150, n149, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(265)
    nor (n2504, n153, n152, byte_counter[5], n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(266)
    nor (n2510, n153, n152, byte_counter[5], n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(267)
    nor (n2516, n153, n152, byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(268)
    nor (n2521, n153, n152, byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(269)
    nor (n2527, n153, n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(270)
    nor (n2532, n153, n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(271)
    nor (n2537, n153, n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(272)
    nor (n2541, n153, n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(273)
    nor (n2548, n153, n152, byte_counter[5], byte_counter[4], n149, 
        n148, n147, n146) ;   // modexp_top.v(274)
    nor (n2554, n153, n152, byte_counter[5], byte_counter[4], n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(275)
    nor (n2560, n153, n152, byte_counter[5], byte_counter[4], n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(276)
    nor (n2565, n153, n152, byte_counter[5], byte_counter[4], n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(277)
    nor (n2571, n153, n152, byte_counter[5], byte_counter[4], n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(278)
    nor (n2576, n153, n152, byte_counter[5], byte_counter[4], n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(279)
    nor (n2581, n153, n152, byte_counter[5], byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(280)
    nor (n2585, n153, n152, byte_counter[5], byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(281)
    nor (n2591, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(282)
    nor (n2596, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(283)
    nor (n2601, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(284)
    nor (n2605, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(285)
    nor (n2610, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(286)
    nor (n2614, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(287)
    nor (n2618, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(288)
    nor (n2621, n153, n152, byte_counter[5], byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(289)
    nor (n2629, n153, byte_counter[6], n151, n150, n149, n148, 
        n147, n146) ;   // modexp_top.v(290)
    nor (n2636, n153, byte_counter[6], n151, n150, n149, n148, 
        n147, byte_counter[0]) ;   // modexp_top.v(291)
    nor (n2643, n153, byte_counter[6], n151, n150, n149, n148, 
        byte_counter[1], n146) ;   // modexp_top.v(292)
    nor (n2649, n153, byte_counter[6], n151, n150, n149, n148, 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(293)
    nor (n2656, n153, byte_counter[6], n151, n150, n149, byte_counter[2], 
        n147, n146) ;   // modexp_top.v(294)
    nor (n2662, n153, byte_counter[6], n151, n150, n149, byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(295)
    nor (n2668, n153, byte_counter[6], n151, n150, n149, byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(296)
    nor (n2673, n153, byte_counter[6], n151, n150, n149, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(297)
    nor (n2680, n153, byte_counter[6], n151, n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(298)
    nor (n2686, n153, byte_counter[6], n151, n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(299)
    nor (n2692, n153, byte_counter[6], n151, n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(300)
    nor (n2697, n153, byte_counter[6], n151, n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(301)
    nor (n2703, n153, byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(302)
    nor (n2708, n153, byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(303)
    nor (n2713, n153, byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(304)
    nor (n2717, n153, byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(305)
    nor (n2724, n153, byte_counter[6], n151, byte_counter[4], n149, 
        n148, n147, n146) ;   // modexp_top.v(306)
    nor (n2730, n153, byte_counter[6], n151, byte_counter[4], n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(307)
    nor (n2736, n153, byte_counter[6], n151, byte_counter[4], n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(308)
    nor (n2741, n153, byte_counter[6], n151, byte_counter[4], n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(309)
    nor (n2747, n153, byte_counter[6], n151, byte_counter[4], n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(310)
    nor (n2752, n153, byte_counter[6], n151, byte_counter[4], n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(311)
    nor (n2757, n153, byte_counter[6], n151, byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(312)
    nor (n2761, n153, byte_counter[6], n151, byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(313)
    nor (n2767, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(314)
    nor (n2772, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(315)
    nor (n2777, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(316)
    nor (n2781, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(317)
    nor (n2786, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(318)
    nor (n2790, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(319)
    nor (n2794, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(320)
    nor (n2797, n153, byte_counter[6], n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(321)
    nor (n2804, n153, byte_counter[6], byte_counter[5], n150, n149, 
        n148, n147, n146) ;   // modexp_top.v(322)
    nor (n2810, n153, byte_counter[6], byte_counter[5], n150, n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(323)
    nor (n2816, n153, byte_counter[6], byte_counter[5], n150, n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(324)
    nor (n2821, n153, byte_counter[6], byte_counter[5], n150, n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(325)
    nor (n2827, n153, byte_counter[6], byte_counter[5], n150, n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(326)
    nor (n2832, n153, byte_counter[6], byte_counter[5], n150, n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(327)
    nor (n2837, n153, byte_counter[6], byte_counter[5], n150, n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(328)
    nor (n2841, n153, byte_counter[6], byte_counter[5], n150, n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(329)
    nor (n2847, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(330)
    nor (n2852, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(331)
    nor (n2857, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(332)
    nor (n2861, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(333)
    nor (n2866, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(334)
    nor (n2870, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(335)
    nor (n2874, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(336)
    nor (n2877, n153, byte_counter[6], byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(337)
    nor (n2883, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, n147, n146) ;   // modexp_top.v(338)
    nor (n2888, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(339)
    nor (n2893, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], n146) ;   // modexp_top.v(340)
    nor (n2897, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(341)
    nor (n2902, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, n146) ;   // modexp_top.v(342)
    nor (n2906, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(343)
    nor (n2910, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(344)
    nor (n2913, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(345)
    nor (n2918, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, n146) ;   // modexp_top.v(346)
    nor (n2922, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, byte_counter[0]) ;   // modexp_top.v(347)
    nor (n2926, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], n146) ;   // modexp_top.v(348)
    nor (n2929, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(349)
    nor (n2933, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, n146) ;   // modexp_top.v(350)
    nor (n2936, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(351)
    nor (n2939, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(352)
    nor (n2941, n153, byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(353)
    nor (n2949, byte_counter[7], n152, n151, n150, n149, n148, 
        n147, n146) ;   // modexp_top.v(354)
    nor (n2956, byte_counter[7], n152, n151, n150, n149, n148, 
        n147, byte_counter[0]) ;   // modexp_top.v(355)
    nor (n2963, byte_counter[7], n152, n151, n150, n149, n148, 
        byte_counter[1], n146) ;   // modexp_top.v(356)
    nor (n2969, byte_counter[7], n152, n151, n150, n149, n148, 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(357)
    nor (n2976, byte_counter[7], n152, n151, n150, n149, byte_counter[2], 
        n147, n146) ;   // modexp_top.v(358)
    nor (n2982, byte_counter[7], n152, n151, n150, n149, byte_counter[2], 
        n147, byte_counter[0]) ;   // modexp_top.v(359)
    nor (n2988, byte_counter[7], n152, n151, n150, n149, byte_counter[2], 
        byte_counter[1], n146) ;   // modexp_top.v(360)
    nor (n2993, byte_counter[7], n152, n151, n150, n149, byte_counter[2], 
        byte_counter[1], byte_counter[0]) ;   // modexp_top.v(361)
    nor (n3000, byte_counter[7], n152, n151, n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(362)
    nor (n3006, byte_counter[7], n152, n151, n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(363)
    nor (n3012, byte_counter[7], n152, n151, n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(364)
    nor (n3017, byte_counter[7], n152, n151, n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(365)
    nor (n3023, byte_counter[7], n152, n151, n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(366)
    nor (n3028, byte_counter[7], n152, n151, n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(367)
    nor (n3033, byte_counter[7], n152, n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(368)
    nor (n3037, byte_counter[7], n152, n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(369)
    nor (n3044, byte_counter[7], n152, n151, byte_counter[4], n149, 
        n148, n147, n146) ;   // modexp_top.v(370)
    nor (n3050, byte_counter[7], n152, n151, byte_counter[4], n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(371)
    nor (n3056, byte_counter[7], n152, n151, byte_counter[4], n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(372)
    nor (n3061, byte_counter[7], n152, n151, byte_counter[4], n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(373)
    nor (n3067, byte_counter[7], n152, n151, byte_counter[4], n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(374)
    nor (n3072, byte_counter[7], n152, n151, byte_counter[4], n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(375)
    nor (n3077, byte_counter[7], n152, n151, byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(376)
    nor (n3081, byte_counter[7], n152, n151, byte_counter[4], n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(377)
    nor (n3087, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(378)
    nor (n3092, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(379)
    nor (n3097, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(380)
    nor (n3101, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(381)
    nor (n3106, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(382)
    nor (n3110, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(383)
    nor (n3114, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(384)
    nor (n3117, byte_counter[7], n152, n151, byte_counter[4], byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(385)
    nor (n3124, byte_counter[7], n152, byte_counter[5], n150, n149, 
        n148, n147, n146) ;   // modexp_top.v(386)
    nor (n3130, byte_counter[7], n152, byte_counter[5], n150, n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(387)
    nor (n3136, byte_counter[7], n152, byte_counter[5], n150, n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(388)
    nor (n3141, byte_counter[7], n152, byte_counter[5], n150, n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(389)
    nor (n3147, byte_counter[7], n152, byte_counter[5], n150, n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(390)
    nor (n3152, byte_counter[7], n152, byte_counter[5], n150, n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(391)
    nor (n3157, byte_counter[7], n152, byte_counter[5], n150, n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(392)
    nor (n3161, byte_counter[7], n152, byte_counter[5], n150, n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(393)
    nor (n3167, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(394)
    nor (n3172, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(395)
    nor (n3177, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(396)
    nor (n3181, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(397)
    nor (n3186, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(398)
    nor (n3190, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(399)
    nor (n3194, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(400)
    nor (n3197, byte_counter[7], n152, byte_counter[5], n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(401)
    nor (n3203, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, n148, n147, n146) ;   // modexp_top.v(402)
    nor (n3208, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(403)
    nor (n3213, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], n146) ;   // modexp_top.v(404)
    nor (n3217, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(405)
    nor (n3222, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, n146) ;   // modexp_top.v(406)
    nor (n3226, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(407)
    nor (n3230, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(408)
    nor (n3233, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(409)
    nor (n3238, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, n146) ;   // modexp_top.v(410)
    nor (n3242, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, byte_counter[0]) ;   // modexp_top.v(411)
    nor (n3246, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], n146) ;   // modexp_top.v(412)
    nor (n3249, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(413)
    nor (n3253, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, n146) ;   // modexp_top.v(414)
    nor (n3256, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(415)
    nor (n3259, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(416)
    nor (n3261, byte_counter[7], n152, byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(417)
    nor (n3268, byte_counter[7], byte_counter[6], n151, n150, n149, 
        n148, n147, n146) ;   // modexp_top.v(418)
    nor (n3274, byte_counter[7], byte_counter[6], n151, n150, n149, 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(419)
    nor (n3280, byte_counter[7], byte_counter[6], n151, n150, n149, 
        n148, byte_counter[1], n146) ;   // modexp_top.v(420)
    nor (n3285, byte_counter[7], byte_counter[6], n151, n150, n149, 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(421)
    nor (n3291, byte_counter[7], byte_counter[6], n151, n150, n149, 
        byte_counter[2], n147, n146) ;   // modexp_top.v(422)
    nor (n3296, byte_counter[7], byte_counter[6], n151, n150, n149, 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(423)
    nor (n3301, byte_counter[7], byte_counter[6], n151, n150, n149, 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(424)
    nor (n3305, byte_counter[7], byte_counter[6], n151, n150, n149, 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(425)
    nor (n3311, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        n148, n147, n146) ;   // modexp_top.v(426)
    nor (n3316, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        n148, n147, byte_counter[0]) ;   // modexp_top.v(427)
    nor (n3321, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        n148, byte_counter[1], n146) ;   // modexp_top.v(428)
    nor (n3325, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(429)
    nor (n3330, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], n147, n146) ;   // modexp_top.v(430)
    nor (n3334, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(431)
    nor (n3338, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(432)
    nor (n3341, byte_counter[7], byte_counter[6], n151, n150, byte_counter[3], 
        byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(433)
    nor (n3347, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, n148, n147, n146) ;   // modexp_top.v(434)
    nor (n3352, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(435)
    nor (n3357, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, n148, byte_counter[1], n146) ;   // modexp_top.v(436)
    nor (n3361, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(437)
    nor (n3366, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, byte_counter[2], n147, n146) ;   // modexp_top.v(438)
    nor (n3370, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(439)
    nor (n3374, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(440)
    nor (n3377, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(441)
    nor (n3382, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], n148, n147, n146) ;   // modexp_top.v(442)
    nor (n3386, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], n148, n147, byte_counter[0]) ;   // modexp_top.v(443)
    nor (n3390, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], n146) ;   // modexp_top.v(444)
    nor (n3393, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(445)
    nor (n3397, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, n146) ;   // modexp_top.v(446)
    nor (n3400, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(447)
    nor (n3403, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(448)
    nor (n3405, byte_counter[7], byte_counter[6], n151, byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(449)
    nor (n3411, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, n148, n147, n146) ;   // modexp_top.v(450)
    nor (n3416, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(451)
    nor (n3421, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, n148, byte_counter[1], n146) ;   // modexp_top.v(452)
    nor (n3425, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(453)
    nor (n3430, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, byte_counter[2], n147, n146) ;   // modexp_top.v(454)
    nor (n3434, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(455)
    nor (n3438, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(456)
    nor (n3441, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        n149, byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(457)
    nor (n3446, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], n148, n147, n146) ;   // modexp_top.v(458)
    nor (n3450, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], n148, n147, byte_counter[0]) ;   // modexp_top.v(459)
    nor (n3454, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], n148, byte_counter[1], n146) ;   // modexp_top.v(460)
    nor (n3457, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(461)
    nor (n3461, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], byte_counter[2], n147, n146) ;   // modexp_top.v(462)
    nor (n3464, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(463)
    nor (n3467, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(464)
    nor (n3469, byte_counter[7], byte_counter[6], byte_counter[5], n150, 
        byte_counter[3], byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(465)
    nor (n3474, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, n147, n146) ;   // modexp_top.v(466)
    nor (n3478, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, n147, byte_counter[0]) ;   // modexp_top.v(467)
    nor (n3482, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], n146) ;   // modexp_top.v(468)
    nor (n3485, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(469)
    nor (n3489, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, n146) ;   // modexp_top.v(470)
    nor (n3492, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(471)
    nor (n3495, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(472)
    nor (n3497, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        n149, byte_counter[2], byte_counter[1], byte_counter[0]) ;   // modexp_top.v(473)
    nor (n3501, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, n146) ;   // modexp_top.v(474)
    nor (n3504, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, n147, byte_counter[0]) ;   // modexp_top.v(475)
    nor (n3507, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], n146) ;   // modexp_top.v(476)
    nor (n3509, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], n148, byte_counter[1], byte_counter[0]) ;   // modexp_top.v(477)
    nor (n3512, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, n146) ;   // modexp_top.v(478)
    nor (n3514, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], n147, byte_counter[0]) ;   // modexp_top.v(479)
    nor (n3516, byte_counter[7], byte_counter[6], byte_counter[5], byte_counter[4], 
        byte_counter[3], byte_counter[2], byte_counter[1], n146) ;   // modexp_top.v(480)
    assign n3517 = n3516 ? encrypted_data_buf[2039] : encrypted_data_buf[2047];   // modexp_top.v(481)
    assign n3518 = n3516 ? encrypted_data_buf[2038] : encrypted_data_buf[2046];   // modexp_top.v(481)
    assign n3519 = n3516 ? encrypted_data_buf[2037] : encrypted_data_buf[2045];   // modexp_top.v(481)
    assign n3520 = n3516 ? encrypted_data_buf[2036] : encrypted_data_buf[2044];   // modexp_top.v(481)
    assign n3521 = n3516 ? encrypted_data_buf[2035] : encrypted_data_buf[2043];   // modexp_top.v(481)
    assign n3522 = n3516 ? encrypted_data_buf[2034] : encrypted_data_buf[2042];   // modexp_top.v(481)
    assign n3523 = n3516 ? encrypted_data_buf[2033] : encrypted_data_buf[2041];   // modexp_top.v(481)
    assign n3524 = n3516 ? encrypted_data_buf[2032] : encrypted_data_buf[2040];   // modexp_top.v(481)
    assign n3525 = n3514 ? encrypted_data_buf[2031] : n3517;   // modexp_top.v(481)
    assign n3526 = n3514 ? encrypted_data_buf[2030] : n3518;   // modexp_top.v(481)
    assign n3527 = n3514 ? encrypted_data_buf[2029] : n3519;   // modexp_top.v(481)
    assign n3528 = n3514 ? encrypted_data_buf[2028] : n3520;   // modexp_top.v(481)
    assign n3529 = n3514 ? encrypted_data_buf[2027] : n3521;   // modexp_top.v(481)
    assign n3530 = n3514 ? encrypted_data_buf[2026] : n3522;   // modexp_top.v(481)
    assign n3531 = n3514 ? encrypted_data_buf[2025] : n3523;   // modexp_top.v(481)
    assign n3532 = n3514 ? encrypted_data_buf[2024] : n3524;   // modexp_top.v(481)
    assign n3533 = n3512 ? encrypted_data_buf[2023] : n3525;   // modexp_top.v(481)
    assign n3534 = n3512 ? encrypted_data_buf[2022] : n3526;   // modexp_top.v(481)
    assign n3535 = n3512 ? encrypted_data_buf[2021] : n3527;   // modexp_top.v(481)
    assign n3536 = n3512 ? encrypted_data_buf[2020] : n3528;   // modexp_top.v(481)
    assign n3537 = n3512 ? encrypted_data_buf[2019] : n3529;   // modexp_top.v(481)
    assign n3538 = n3512 ? encrypted_data_buf[2018] : n3530;   // modexp_top.v(481)
    assign n3539 = n3512 ? encrypted_data_buf[2017] : n3531;   // modexp_top.v(481)
    assign n3540 = n3512 ? encrypted_data_buf[2016] : n3532;   // modexp_top.v(481)
    assign n3541 = n3509 ? encrypted_data_buf[2015] : n3533;   // modexp_top.v(481)
    assign n3542 = n3509 ? encrypted_data_buf[2014] : n3534;   // modexp_top.v(481)
    assign n3543 = n3509 ? encrypted_data_buf[2013] : n3535;   // modexp_top.v(481)
    assign n3544 = n3509 ? encrypted_data_buf[2012] : n3536;   // modexp_top.v(481)
    assign n3545 = n3509 ? encrypted_data_buf[2011] : n3537;   // modexp_top.v(481)
    assign n3546 = n3509 ? encrypted_data_buf[2010] : n3538;   // modexp_top.v(481)
    assign n3547 = n3509 ? encrypted_data_buf[2009] : n3539;   // modexp_top.v(481)
    assign n3548 = n3509 ? encrypted_data_buf[2008] : n3540;   // modexp_top.v(481)
    assign n3549 = n3507 ? encrypted_data_buf[2007] : n3541;   // modexp_top.v(481)
    assign n3550 = n3507 ? encrypted_data_buf[2006] : n3542;   // modexp_top.v(481)
    assign n3551 = n3507 ? encrypted_data_buf[2005] : n3543;   // modexp_top.v(481)
    assign n3552 = n3507 ? encrypted_data_buf[2004] : n3544;   // modexp_top.v(481)
    assign n3553 = n3507 ? encrypted_data_buf[2003] : n3545;   // modexp_top.v(481)
    assign n3554 = n3507 ? encrypted_data_buf[2002] : n3546;   // modexp_top.v(481)
    assign n3555 = n3507 ? encrypted_data_buf[2001] : n3547;   // modexp_top.v(481)
    assign n3556 = n3507 ? encrypted_data_buf[2000] : n3548;   // modexp_top.v(481)
    assign n3557 = n3504 ? encrypted_data_buf[1999] : n3549;   // modexp_top.v(481)
    assign n3558 = n3504 ? encrypted_data_buf[1998] : n3550;   // modexp_top.v(481)
    assign n3559 = n3504 ? encrypted_data_buf[1997] : n3551;   // modexp_top.v(481)
    assign n3560 = n3504 ? encrypted_data_buf[1996] : n3552;   // modexp_top.v(481)
    assign n3561 = n3504 ? encrypted_data_buf[1995] : n3553;   // modexp_top.v(481)
    assign n3562 = n3504 ? encrypted_data_buf[1994] : n3554;   // modexp_top.v(481)
    assign n3563 = n3504 ? encrypted_data_buf[1993] : n3555;   // modexp_top.v(481)
    assign n3564 = n3504 ? encrypted_data_buf[1992] : n3556;   // modexp_top.v(481)
    assign n3565 = n3501 ? encrypted_data_buf[1991] : n3557;   // modexp_top.v(481)
    assign n3566 = n3501 ? encrypted_data_buf[1990] : n3558;   // modexp_top.v(481)
    assign n3567 = n3501 ? encrypted_data_buf[1989] : n3559;   // modexp_top.v(481)
    assign n3568 = n3501 ? encrypted_data_buf[1988] : n3560;   // modexp_top.v(481)
    assign n3569 = n3501 ? encrypted_data_buf[1987] : n3561;   // modexp_top.v(481)
    assign n3570 = n3501 ? encrypted_data_buf[1986] : n3562;   // modexp_top.v(481)
    assign n3571 = n3501 ? encrypted_data_buf[1985] : n3563;   // modexp_top.v(481)
    assign n3572 = n3501 ? encrypted_data_buf[1984] : n3564;   // modexp_top.v(481)
    assign n3573 = n3497 ? encrypted_data_buf[1983] : n3565;   // modexp_top.v(481)
    assign n3574 = n3497 ? encrypted_data_buf[1982] : n3566;   // modexp_top.v(481)
    assign n3575 = n3497 ? encrypted_data_buf[1981] : n3567;   // modexp_top.v(481)
    assign n3576 = n3497 ? encrypted_data_buf[1980] : n3568;   // modexp_top.v(481)
    assign n3577 = n3497 ? encrypted_data_buf[1979] : n3569;   // modexp_top.v(481)
    assign n3578 = n3497 ? encrypted_data_buf[1978] : n3570;   // modexp_top.v(481)
    assign n3579 = n3497 ? encrypted_data_buf[1977] : n3571;   // modexp_top.v(481)
    assign n3580 = n3497 ? encrypted_data_buf[1976] : n3572;   // modexp_top.v(481)
    assign n3581 = n3495 ? encrypted_data_buf[1975] : n3573;   // modexp_top.v(481)
    assign n3582 = n3495 ? encrypted_data_buf[1974] : n3574;   // modexp_top.v(481)
    assign n3583 = n3495 ? encrypted_data_buf[1973] : n3575;   // modexp_top.v(481)
    assign n3584 = n3495 ? encrypted_data_buf[1972] : n3576;   // modexp_top.v(481)
    assign n3585 = n3495 ? encrypted_data_buf[1971] : n3577;   // modexp_top.v(481)
    assign n3586 = n3495 ? encrypted_data_buf[1970] : n3578;   // modexp_top.v(481)
    assign n3587 = n3495 ? encrypted_data_buf[1969] : n3579;   // modexp_top.v(481)
    assign n3588 = n3495 ? encrypted_data_buf[1968] : n3580;   // modexp_top.v(481)
    assign n3589 = n3492 ? encrypted_data_buf[1967] : n3581;   // modexp_top.v(481)
    assign n3590 = n3492 ? encrypted_data_buf[1966] : n3582;   // modexp_top.v(481)
    assign n3591 = n3492 ? encrypted_data_buf[1965] : n3583;   // modexp_top.v(481)
    assign n3592 = n3492 ? encrypted_data_buf[1964] : n3584;   // modexp_top.v(481)
    assign n3593 = n3492 ? encrypted_data_buf[1963] : n3585;   // modexp_top.v(481)
    assign n3594 = n3492 ? encrypted_data_buf[1962] : n3586;   // modexp_top.v(481)
    assign n3595 = n3492 ? encrypted_data_buf[1961] : n3587;   // modexp_top.v(481)
    assign n3596 = n3492 ? encrypted_data_buf[1960] : n3588;   // modexp_top.v(481)
    assign n3597 = n3489 ? encrypted_data_buf[1959] : n3589;   // modexp_top.v(481)
    assign n3598 = n3489 ? encrypted_data_buf[1958] : n3590;   // modexp_top.v(481)
    assign n3599 = n3489 ? encrypted_data_buf[1957] : n3591;   // modexp_top.v(481)
    assign n3600 = n3489 ? encrypted_data_buf[1956] : n3592;   // modexp_top.v(481)
    assign n3601 = n3489 ? encrypted_data_buf[1955] : n3593;   // modexp_top.v(481)
    assign n3602 = n3489 ? encrypted_data_buf[1954] : n3594;   // modexp_top.v(481)
    assign n3603 = n3489 ? encrypted_data_buf[1953] : n3595;   // modexp_top.v(481)
    assign n3604 = n3489 ? encrypted_data_buf[1952] : n3596;   // modexp_top.v(481)
    assign n3605 = n3485 ? encrypted_data_buf[1951] : n3597;   // modexp_top.v(481)
    assign n3606 = n3485 ? encrypted_data_buf[1950] : n3598;   // modexp_top.v(481)
    assign n3607 = n3485 ? encrypted_data_buf[1949] : n3599;   // modexp_top.v(481)
    assign n3608 = n3485 ? encrypted_data_buf[1948] : n3600;   // modexp_top.v(481)
    assign n3609 = n3485 ? encrypted_data_buf[1947] : n3601;   // modexp_top.v(481)
    assign n3610 = n3485 ? encrypted_data_buf[1946] : n3602;   // modexp_top.v(481)
    assign n3611 = n3485 ? encrypted_data_buf[1945] : n3603;   // modexp_top.v(481)
    assign n3612 = n3485 ? encrypted_data_buf[1944] : n3604;   // modexp_top.v(481)
    assign n3613 = n3482 ? encrypted_data_buf[1943] : n3605;   // modexp_top.v(481)
    assign n3614 = n3482 ? encrypted_data_buf[1942] : n3606;   // modexp_top.v(481)
    assign n3615 = n3482 ? encrypted_data_buf[1941] : n3607;   // modexp_top.v(481)
    assign n3616 = n3482 ? encrypted_data_buf[1940] : n3608;   // modexp_top.v(481)
    assign n3617 = n3482 ? encrypted_data_buf[1939] : n3609;   // modexp_top.v(481)
    assign n3618 = n3482 ? encrypted_data_buf[1938] : n3610;   // modexp_top.v(481)
    assign n3619 = n3482 ? encrypted_data_buf[1937] : n3611;   // modexp_top.v(481)
    assign n3620 = n3482 ? encrypted_data_buf[1936] : n3612;   // modexp_top.v(481)
    assign n3621 = n3478 ? encrypted_data_buf[1935] : n3613;   // modexp_top.v(481)
    assign n3622 = n3478 ? encrypted_data_buf[1934] : n3614;   // modexp_top.v(481)
    assign n3623 = n3478 ? encrypted_data_buf[1933] : n3615;   // modexp_top.v(481)
    assign n3624 = n3478 ? encrypted_data_buf[1932] : n3616;   // modexp_top.v(481)
    assign n3625 = n3478 ? encrypted_data_buf[1931] : n3617;   // modexp_top.v(481)
    assign n3626 = n3478 ? encrypted_data_buf[1930] : n3618;   // modexp_top.v(481)
    assign n3627 = n3478 ? encrypted_data_buf[1929] : n3619;   // modexp_top.v(481)
    assign n3628 = n3478 ? encrypted_data_buf[1928] : n3620;   // modexp_top.v(481)
    assign n3629 = n3474 ? encrypted_data_buf[1927] : n3621;   // modexp_top.v(481)
    assign n3630 = n3474 ? encrypted_data_buf[1926] : n3622;   // modexp_top.v(481)
    assign n3631 = n3474 ? encrypted_data_buf[1925] : n3623;   // modexp_top.v(481)
    assign n3632 = n3474 ? encrypted_data_buf[1924] : n3624;   // modexp_top.v(481)
    assign n3633 = n3474 ? encrypted_data_buf[1923] : n3625;   // modexp_top.v(481)
    assign n3634 = n3474 ? encrypted_data_buf[1922] : n3626;   // modexp_top.v(481)
    assign n3635 = n3474 ? encrypted_data_buf[1921] : n3627;   // modexp_top.v(481)
    assign n3636 = n3474 ? encrypted_data_buf[1920] : n3628;   // modexp_top.v(481)
    assign n3637 = n3469 ? encrypted_data_buf[1919] : n3629;   // modexp_top.v(481)
    assign n3638 = n3469 ? encrypted_data_buf[1918] : n3630;   // modexp_top.v(481)
    assign n3639 = n3469 ? encrypted_data_buf[1917] : n3631;   // modexp_top.v(481)
    assign n3640 = n3469 ? encrypted_data_buf[1916] : n3632;   // modexp_top.v(481)
    assign n3641 = n3469 ? encrypted_data_buf[1915] : n3633;   // modexp_top.v(481)
    assign n3642 = n3469 ? encrypted_data_buf[1914] : n3634;   // modexp_top.v(481)
    assign n3643 = n3469 ? encrypted_data_buf[1913] : n3635;   // modexp_top.v(481)
    assign n3644 = n3469 ? encrypted_data_buf[1912] : n3636;   // modexp_top.v(481)
    assign n3645 = n3467 ? encrypted_data_buf[1911] : n3637;   // modexp_top.v(481)
    assign n3646 = n3467 ? encrypted_data_buf[1910] : n3638;   // modexp_top.v(481)
    assign n3647 = n3467 ? encrypted_data_buf[1909] : n3639;   // modexp_top.v(481)
    assign n3648 = n3467 ? encrypted_data_buf[1908] : n3640;   // modexp_top.v(481)
    assign n3649 = n3467 ? encrypted_data_buf[1907] : n3641;   // modexp_top.v(481)
    assign n3650 = n3467 ? encrypted_data_buf[1906] : n3642;   // modexp_top.v(481)
    assign n3651 = n3467 ? encrypted_data_buf[1905] : n3643;   // modexp_top.v(481)
    assign n3652 = n3467 ? encrypted_data_buf[1904] : n3644;   // modexp_top.v(481)
    assign n3653 = n3464 ? encrypted_data_buf[1903] : n3645;   // modexp_top.v(481)
    assign n3654 = n3464 ? encrypted_data_buf[1902] : n3646;   // modexp_top.v(481)
    assign n3655 = n3464 ? encrypted_data_buf[1901] : n3647;   // modexp_top.v(481)
    assign n3656 = n3464 ? encrypted_data_buf[1900] : n3648;   // modexp_top.v(481)
    assign n3657 = n3464 ? encrypted_data_buf[1899] : n3649;   // modexp_top.v(481)
    assign n3658 = n3464 ? encrypted_data_buf[1898] : n3650;   // modexp_top.v(481)
    assign n3659 = n3464 ? encrypted_data_buf[1897] : n3651;   // modexp_top.v(481)
    assign n3660 = n3464 ? encrypted_data_buf[1896] : n3652;   // modexp_top.v(481)
    assign n3661 = n3461 ? encrypted_data_buf[1895] : n3653;   // modexp_top.v(481)
    assign n3662 = n3461 ? encrypted_data_buf[1894] : n3654;   // modexp_top.v(481)
    assign n3663 = n3461 ? encrypted_data_buf[1893] : n3655;   // modexp_top.v(481)
    assign n3664 = n3461 ? encrypted_data_buf[1892] : n3656;   // modexp_top.v(481)
    assign n3665 = n3461 ? encrypted_data_buf[1891] : n3657;   // modexp_top.v(481)
    assign n3666 = n3461 ? encrypted_data_buf[1890] : n3658;   // modexp_top.v(481)
    assign n3667 = n3461 ? encrypted_data_buf[1889] : n3659;   // modexp_top.v(481)
    assign n3668 = n3461 ? encrypted_data_buf[1888] : n3660;   // modexp_top.v(481)
    assign n3669 = n3457 ? encrypted_data_buf[1887] : n3661;   // modexp_top.v(481)
    assign n3670 = n3457 ? encrypted_data_buf[1886] : n3662;   // modexp_top.v(481)
    assign n3671 = n3457 ? encrypted_data_buf[1885] : n3663;   // modexp_top.v(481)
    assign n3672 = n3457 ? encrypted_data_buf[1884] : n3664;   // modexp_top.v(481)
    assign n3673 = n3457 ? encrypted_data_buf[1883] : n3665;   // modexp_top.v(481)
    assign n3674 = n3457 ? encrypted_data_buf[1882] : n3666;   // modexp_top.v(481)
    assign n3675 = n3457 ? encrypted_data_buf[1881] : n3667;   // modexp_top.v(481)
    assign n3676 = n3457 ? encrypted_data_buf[1880] : n3668;   // modexp_top.v(481)
    assign n3677 = n3454 ? encrypted_data_buf[1879] : n3669;   // modexp_top.v(481)
    assign n3678 = n3454 ? encrypted_data_buf[1878] : n3670;   // modexp_top.v(481)
    assign n3679 = n3454 ? encrypted_data_buf[1877] : n3671;   // modexp_top.v(481)
    assign n3680 = n3454 ? encrypted_data_buf[1876] : n3672;   // modexp_top.v(481)
    assign n3681 = n3454 ? encrypted_data_buf[1875] : n3673;   // modexp_top.v(481)
    assign n3682 = n3454 ? encrypted_data_buf[1874] : n3674;   // modexp_top.v(481)
    assign n3683 = n3454 ? encrypted_data_buf[1873] : n3675;   // modexp_top.v(481)
    assign n3684 = n3454 ? encrypted_data_buf[1872] : n3676;   // modexp_top.v(481)
    assign n3685 = n3450 ? encrypted_data_buf[1871] : n3677;   // modexp_top.v(481)
    assign n3686 = n3450 ? encrypted_data_buf[1870] : n3678;   // modexp_top.v(481)
    assign n3687 = n3450 ? encrypted_data_buf[1869] : n3679;   // modexp_top.v(481)
    assign n3688 = n3450 ? encrypted_data_buf[1868] : n3680;   // modexp_top.v(481)
    assign n3689 = n3450 ? encrypted_data_buf[1867] : n3681;   // modexp_top.v(481)
    assign n3690 = n3450 ? encrypted_data_buf[1866] : n3682;   // modexp_top.v(481)
    assign n3691 = n3450 ? encrypted_data_buf[1865] : n3683;   // modexp_top.v(481)
    assign n3692 = n3450 ? encrypted_data_buf[1864] : n3684;   // modexp_top.v(481)
    assign n3693 = n3446 ? encrypted_data_buf[1863] : n3685;   // modexp_top.v(481)
    assign n3694 = n3446 ? encrypted_data_buf[1862] : n3686;   // modexp_top.v(481)
    assign n3695 = n3446 ? encrypted_data_buf[1861] : n3687;   // modexp_top.v(481)
    assign n3696 = n3446 ? encrypted_data_buf[1860] : n3688;   // modexp_top.v(481)
    assign n3697 = n3446 ? encrypted_data_buf[1859] : n3689;   // modexp_top.v(481)
    assign n3698 = n3446 ? encrypted_data_buf[1858] : n3690;   // modexp_top.v(481)
    assign n3699 = n3446 ? encrypted_data_buf[1857] : n3691;   // modexp_top.v(481)
    assign n3700 = n3446 ? encrypted_data_buf[1856] : n3692;   // modexp_top.v(481)
    assign n3701 = n3441 ? encrypted_data_buf[1855] : n3693;   // modexp_top.v(481)
    assign n3702 = n3441 ? encrypted_data_buf[1854] : n3694;   // modexp_top.v(481)
    assign n3703 = n3441 ? encrypted_data_buf[1853] : n3695;   // modexp_top.v(481)
    assign n3704 = n3441 ? encrypted_data_buf[1852] : n3696;   // modexp_top.v(481)
    assign n3705 = n3441 ? encrypted_data_buf[1851] : n3697;   // modexp_top.v(481)
    assign n3706 = n3441 ? encrypted_data_buf[1850] : n3698;   // modexp_top.v(481)
    assign n3707 = n3441 ? encrypted_data_buf[1849] : n3699;   // modexp_top.v(481)
    assign n3708 = n3441 ? encrypted_data_buf[1848] : n3700;   // modexp_top.v(481)
    assign n3709 = n3438 ? encrypted_data_buf[1847] : n3701;   // modexp_top.v(481)
    assign n3710 = n3438 ? encrypted_data_buf[1846] : n3702;   // modexp_top.v(481)
    assign n3711 = n3438 ? encrypted_data_buf[1845] : n3703;   // modexp_top.v(481)
    assign n3712 = n3438 ? encrypted_data_buf[1844] : n3704;   // modexp_top.v(481)
    assign n3713 = n3438 ? encrypted_data_buf[1843] : n3705;   // modexp_top.v(481)
    assign n3714 = n3438 ? encrypted_data_buf[1842] : n3706;   // modexp_top.v(481)
    assign n3715 = n3438 ? encrypted_data_buf[1841] : n3707;   // modexp_top.v(481)
    assign n3716 = n3438 ? encrypted_data_buf[1840] : n3708;   // modexp_top.v(481)
    assign n3717 = n3434 ? encrypted_data_buf[1839] : n3709;   // modexp_top.v(481)
    assign n3718 = n3434 ? encrypted_data_buf[1838] : n3710;   // modexp_top.v(481)
    assign n3719 = n3434 ? encrypted_data_buf[1837] : n3711;   // modexp_top.v(481)
    assign n3720 = n3434 ? encrypted_data_buf[1836] : n3712;   // modexp_top.v(481)
    assign n3721 = n3434 ? encrypted_data_buf[1835] : n3713;   // modexp_top.v(481)
    assign n3722 = n3434 ? encrypted_data_buf[1834] : n3714;   // modexp_top.v(481)
    assign n3723 = n3434 ? encrypted_data_buf[1833] : n3715;   // modexp_top.v(481)
    assign n3724 = n3434 ? encrypted_data_buf[1832] : n3716;   // modexp_top.v(481)
    assign n3725 = n3430 ? encrypted_data_buf[1831] : n3717;   // modexp_top.v(481)
    assign n3726 = n3430 ? encrypted_data_buf[1830] : n3718;   // modexp_top.v(481)
    assign n3727 = n3430 ? encrypted_data_buf[1829] : n3719;   // modexp_top.v(481)
    assign n3728 = n3430 ? encrypted_data_buf[1828] : n3720;   // modexp_top.v(481)
    assign n3729 = n3430 ? encrypted_data_buf[1827] : n3721;   // modexp_top.v(481)
    assign n3730 = n3430 ? encrypted_data_buf[1826] : n3722;   // modexp_top.v(481)
    assign n3731 = n3430 ? encrypted_data_buf[1825] : n3723;   // modexp_top.v(481)
    assign n3732 = n3430 ? encrypted_data_buf[1824] : n3724;   // modexp_top.v(481)
    assign n3733 = n3425 ? encrypted_data_buf[1823] : n3725;   // modexp_top.v(481)
    assign n3734 = n3425 ? encrypted_data_buf[1822] : n3726;   // modexp_top.v(481)
    assign n3735 = n3425 ? encrypted_data_buf[1821] : n3727;   // modexp_top.v(481)
    assign n3736 = n3425 ? encrypted_data_buf[1820] : n3728;   // modexp_top.v(481)
    assign n3737 = n3425 ? encrypted_data_buf[1819] : n3729;   // modexp_top.v(481)
    assign n3738 = n3425 ? encrypted_data_buf[1818] : n3730;   // modexp_top.v(481)
    assign n3739 = n3425 ? encrypted_data_buf[1817] : n3731;   // modexp_top.v(481)
    assign n3740 = n3425 ? encrypted_data_buf[1816] : n3732;   // modexp_top.v(481)
    assign n3741 = n3421 ? encrypted_data_buf[1815] : n3733;   // modexp_top.v(481)
    assign n3742 = n3421 ? encrypted_data_buf[1814] : n3734;   // modexp_top.v(481)
    assign n3743 = n3421 ? encrypted_data_buf[1813] : n3735;   // modexp_top.v(481)
    assign n3744 = n3421 ? encrypted_data_buf[1812] : n3736;   // modexp_top.v(481)
    assign n3745 = n3421 ? encrypted_data_buf[1811] : n3737;   // modexp_top.v(481)
    assign n3746 = n3421 ? encrypted_data_buf[1810] : n3738;   // modexp_top.v(481)
    assign n3747 = n3421 ? encrypted_data_buf[1809] : n3739;   // modexp_top.v(481)
    assign n3748 = n3421 ? encrypted_data_buf[1808] : n3740;   // modexp_top.v(481)
    assign n3749 = n3416 ? encrypted_data_buf[1807] : n3741;   // modexp_top.v(481)
    assign n3750 = n3416 ? encrypted_data_buf[1806] : n3742;   // modexp_top.v(481)
    assign n3751 = n3416 ? encrypted_data_buf[1805] : n3743;   // modexp_top.v(481)
    assign n3752 = n3416 ? encrypted_data_buf[1804] : n3744;   // modexp_top.v(481)
    assign n3753 = n3416 ? encrypted_data_buf[1803] : n3745;   // modexp_top.v(481)
    assign n3754 = n3416 ? encrypted_data_buf[1802] : n3746;   // modexp_top.v(481)
    assign n3755 = n3416 ? encrypted_data_buf[1801] : n3747;   // modexp_top.v(481)
    assign n3756 = n3416 ? encrypted_data_buf[1800] : n3748;   // modexp_top.v(481)
    assign n3757 = n3411 ? encrypted_data_buf[1799] : n3749;   // modexp_top.v(481)
    assign n3758 = n3411 ? encrypted_data_buf[1798] : n3750;   // modexp_top.v(481)
    assign n3759 = n3411 ? encrypted_data_buf[1797] : n3751;   // modexp_top.v(481)
    assign n3760 = n3411 ? encrypted_data_buf[1796] : n3752;   // modexp_top.v(481)
    assign n3761 = n3411 ? encrypted_data_buf[1795] : n3753;   // modexp_top.v(481)
    assign n3762 = n3411 ? encrypted_data_buf[1794] : n3754;   // modexp_top.v(481)
    assign n3763 = n3411 ? encrypted_data_buf[1793] : n3755;   // modexp_top.v(481)
    assign n3764 = n3411 ? encrypted_data_buf[1792] : n3756;   // modexp_top.v(481)
    assign n3765 = n3405 ? encrypted_data_buf[1791] : n3757;   // modexp_top.v(481)
    assign n3766 = n3405 ? encrypted_data_buf[1790] : n3758;   // modexp_top.v(481)
    assign n3767 = n3405 ? encrypted_data_buf[1789] : n3759;   // modexp_top.v(481)
    assign n3768 = n3405 ? encrypted_data_buf[1788] : n3760;   // modexp_top.v(481)
    assign n3769 = n3405 ? encrypted_data_buf[1787] : n3761;   // modexp_top.v(481)
    assign n3770 = n3405 ? encrypted_data_buf[1786] : n3762;   // modexp_top.v(481)
    assign n3771 = n3405 ? encrypted_data_buf[1785] : n3763;   // modexp_top.v(481)
    assign n3772 = n3405 ? encrypted_data_buf[1784] : n3764;   // modexp_top.v(481)
    assign n3773 = n3403 ? encrypted_data_buf[1783] : n3765;   // modexp_top.v(481)
    assign n3774 = n3403 ? encrypted_data_buf[1782] : n3766;   // modexp_top.v(481)
    assign n3775 = n3403 ? encrypted_data_buf[1781] : n3767;   // modexp_top.v(481)
    assign n3776 = n3403 ? encrypted_data_buf[1780] : n3768;   // modexp_top.v(481)
    assign n3777 = n3403 ? encrypted_data_buf[1779] : n3769;   // modexp_top.v(481)
    assign n3778 = n3403 ? encrypted_data_buf[1778] : n3770;   // modexp_top.v(481)
    assign n3779 = n3403 ? encrypted_data_buf[1777] : n3771;   // modexp_top.v(481)
    assign n3780 = n3403 ? encrypted_data_buf[1776] : n3772;   // modexp_top.v(481)
    assign n3781 = n3400 ? encrypted_data_buf[1775] : n3773;   // modexp_top.v(481)
    assign n3782 = n3400 ? encrypted_data_buf[1774] : n3774;   // modexp_top.v(481)
    assign n3783 = n3400 ? encrypted_data_buf[1773] : n3775;   // modexp_top.v(481)
    assign n3784 = n3400 ? encrypted_data_buf[1772] : n3776;   // modexp_top.v(481)
    assign n3785 = n3400 ? encrypted_data_buf[1771] : n3777;   // modexp_top.v(481)
    assign n3786 = n3400 ? encrypted_data_buf[1770] : n3778;   // modexp_top.v(481)
    assign n3787 = n3400 ? encrypted_data_buf[1769] : n3779;   // modexp_top.v(481)
    assign n3788 = n3400 ? encrypted_data_buf[1768] : n3780;   // modexp_top.v(481)
    assign n3789 = n3397 ? encrypted_data_buf[1767] : n3781;   // modexp_top.v(481)
    assign n3790 = n3397 ? encrypted_data_buf[1766] : n3782;   // modexp_top.v(481)
    assign n3791 = n3397 ? encrypted_data_buf[1765] : n3783;   // modexp_top.v(481)
    assign n3792 = n3397 ? encrypted_data_buf[1764] : n3784;   // modexp_top.v(481)
    assign n3793 = n3397 ? encrypted_data_buf[1763] : n3785;   // modexp_top.v(481)
    assign n3794 = n3397 ? encrypted_data_buf[1762] : n3786;   // modexp_top.v(481)
    assign n3795 = n3397 ? encrypted_data_buf[1761] : n3787;   // modexp_top.v(481)
    assign n3796 = n3397 ? encrypted_data_buf[1760] : n3788;   // modexp_top.v(481)
    assign n3797 = n3393 ? encrypted_data_buf[1759] : n3789;   // modexp_top.v(481)
    assign n3798 = n3393 ? encrypted_data_buf[1758] : n3790;   // modexp_top.v(481)
    assign n3799 = n3393 ? encrypted_data_buf[1757] : n3791;   // modexp_top.v(481)
    assign n3800 = n3393 ? encrypted_data_buf[1756] : n3792;   // modexp_top.v(481)
    assign n3801 = n3393 ? encrypted_data_buf[1755] : n3793;   // modexp_top.v(481)
    assign n3802 = n3393 ? encrypted_data_buf[1754] : n3794;   // modexp_top.v(481)
    assign n3803 = n3393 ? encrypted_data_buf[1753] : n3795;   // modexp_top.v(481)
    assign n3804 = n3393 ? encrypted_data_buf[1752] : n3796;   // modexp_top.v(481)
    assign n3805 = n3390 ? encrypted_data_buf[1751] : n3797;   // modexp_top.v(481)
    assign n3806 = n3390 ? encrypted_data_buf[1750] : n3798;   // modexp_top.v(481)
    assign n3807 = n3390 ? encrypted_data_buf[1749] : n3799;   // modexp_top.v(481)
    assign n3808 = n3390 ? encrypted_data_buf[1748] : n3800;   // modexp_top.v(481)
    assign n3809 = n3390 ? encrypted_data_buf[1747] : n3801;   // modexp_top.v(481)
    assign n3810 = n3390 ? encrypted_data_buf[1746] : n3802;   // modexp_top.v(481)
    assign n3811 = n3390 ? encrypted_data_buf[1745] : n3803;   // modexp_top.v(481)
    assign n3812 = n3390 ? encrypted_data_buf[1744] : n3804;   // modexp_top.v(481)
    assign n3813 = n3386 ? encrypted_data_buf[1743] : n3805;   // modexp_top.v(481)
    assign n3814 = n3386 ? encrypted_data_buf[1742] : n3806;   // modexp_top.v(481)
    assign n3815 = n3386 ? encrypted_data_buf[1741] : n3807;   // modexp_top.v(481)
    assign n3816 = n3386 ? encrypted_data_buf[1740] : n3808;   // modexp_top.v(481)
    assign n3817 = n3386 ? encrypted_data_buf[1739] : n3809;   // modexp_top.v(481)
    assign n3818 = n3386 ? encrypted_data_buf[1738] : n3810;   // modexp_top.v(481)
    assign n3819 = n3386 ? encrypted_data_buf[1737] : n3811;   // modexp_top.v(481)
    assign n3820 = n3386 ? encrypted_data_buf[1736] : n3812;   // modexp_top.v(481)
    assign n3821 = n3382 ? encrypted_data_buf[1735] : n3813;   // modexp_top.v(481)
    assign n3822 = n3382 ? encrypted_data_buf[1734] : n3814;   // modexp_top.v(481)
    assign n3823 = n3382 ? encrypted_data_buf[1733] : n3815;   // modexp_top.v(481)
    assign n3824 = n3382 ? encrypted_data_buf[1732] : n3816;   // modexp_top.v(481)
    assign n3825 = n3382 ? encrypted_data_buf[1731] : n3817;   // modexp_top.v(481)
    assign n3826 = n3382 ? encrypted_data_buf[1730] : n3818;   // modexp_top.v(481)
    assign n3827 = n3382 ? encrypted_data_buf[1729] : n3819;   // modexp_top.v(481)
    assign n3828 = n3382 ? encrypted_data_buf[1728] : n3820;   // modexp_top.v(481)
    assign n3829 = n3377 ? encrypted_data_buf[1727] : n3821;   // modexp_top.v(481)
    assign n3830 = n3377 ? encrypted_data_buf[1726] : n3822;   // modexp_top.v(481)
    assign n3831 = n3377 ? encrypted_data_buf[1725] : n3823;   // modexp_top.v(481)
    assign n3832 = n3377 ? encrypted_data_buf[1724] : n3824;   // modexp_top.v(481)
    assign n3833 = n3377 ? encrypted_data_buf[1723] : n3825;   // modexp_top.v(481)
    assign n3834 = n3377 ? encrypted_data_buf[1722] : n3826;   // modexp_top.v(481)
    assign n3835 = n3377 ? encrypted_data_buf[1721] : n3827;   // modexp_top.v(481)
    assign n3836 = n3377 ? encrypted_data_buf[1720] : n3828;   // modexp_top.v(481)
    assign n3837 = n3374 ? encrypted_data_buf[1719] : n3829;   // modexp_top.v(481)
    assign n3838 = n3374 ? encrypted_data_buf[1718] : n3830;   // modexp_top.v(481)
    assign n3839 = n3374 ? encrypted_data_buf[1717] : n3831;   // modexp_top.v(481)
    assign n3840 = n3374 ? encrypted_data_buf[1716] : n3832;   // modexp_top.v(481)
    assign n3841 = n3374 ? encrypted_data_buf[1715] : n3833;   // modexp_top.v(481)
    assign n3842 = n3374 ? encrypted_data_buf[1714] : n3834;   // modexp_top.v(481)
    assign n3843 = n3374 ? encrypted_data_buf[1713] : n3835;   // modexp_top.v(481)
    assign n3844 = n3374 ? encrypted_data_buf[1712] : n3836;   // modexp_top.v(481)
    assign n3845 = n3370 ? encrypted_data_buf[1711] : n3837;   // modexp_top.v(481)
    assign n3846 = n3370 ? encrypted_data_buf[1710] : n3838;   // modexp_top.v(481)
    assign n3847 = n3370 ? encrypted_data_buf[1709] : n3839;   // modexp_top.v(481)
    assign n3848 = n3370 ? encrypted_data_buf[1708] : n3840;   // modexp_top.v(481)
    assign n3849 = n3370 ? encrypted_data_buf[1707] : n3841;   // modexp_top.v(481)
    assign n3850 = n3370 ? encrypted_data_buf[1706] : n3842;   // modexp_top.v(481)
    assign n3851 = n3370 ? encrypted_data_buf[1705] : n3843;   // modexp_top.v(481)
    assign n3852 = n3370 ? encrypted_data_buf[1704] : n3844;   // modexp_top.v(481)
    assign n3853 = n3366 ? encrypted_data_buf[1703] : n3845;   // modexp_top.v(481)
    assign n3854 = n3366 ? encrypted_data_buf[1702] : n3846;   // modexp_top.v(481)
    assign n3855 = n3366 ? encrypted_data_buf[1701] : n3847;   // modexp_top.v(481)
    assign n3856 = n3366 ? encrypted_data_buf[1700] : n3848;   // modexp_top.v(481)
    assign n3857 = n3366 ? encrypted_data_buf[1699] : n3849;   // modexp_top.v(481)
    assign n3858 = n3366 ? encrypted_data_buf[1698] : n3850;   // modexp_top.v(481)
    assign n3859 = n3366 ? encrypted_data_buf[1697] : n3851;   // modexp_top.v(481)
    assign n3860 = n3366 ? encrypted_data_buf[1696] : n3852;   // modexp_top.v(481)
    assign n3861 = n3361 ? encrypted_data_buf[1695] : n3853;   // modexp_top.v(481)
    assign n3862 = n3361 ? encrypted_data_buf[1694] : n3854;   // modexp_top.v(481)
    assign n3863 = n3361 ? encrypted_data_buf[1693] : n3855;   // modexp_top.v(481)
    assign n3864 = n3361 ? encrypted_data_buf[1692] : n3856;   // modexp_top.v(481)
    assign n3865 = n3361 ? encrypted_data_buf[1691] : n3857;   // modexp_top.v(481)
    assign n3866 = n3361 ? encrypted_data_buf[1690] : n3858;   // modexp_top.v(481)
    assign n3867 = n3361 ? encrypted_data_buf[1689] : n3859;   // modexp_top.v(481)
    assign n3868 = n3361 ? encrypted_data_buf[1688] : n3860;   // modexp_top.v(481)
    assign n3869 = n3357 ? encrypted_data_buf[1687] : n3861;   // modexp_top.v(481)
    assign n3870 = n3357 ? encrypted_data_buf[1686] : n3862;   // modexp_top.v(481)
    assign n3871 = n3357 ? encrypted_data_buf[1685] : n3863;   // modexp_top.v(481)
    assign n3872 = n3357 ? encrypted_data_buf[1684] : n3864;   // modexp_top.v(481)
    assign n3873 = n3357 ? encrypted_data_buf[1683] : n3865;   // modexp_top.v(481)
    assign n3874 = n3357 ? encrypted_data_buf[1682] : n3866;   // modexp_top.v(481)
    assign n3875 = n3357 ? encrypted_data_buf[1681] : n3867;   // modexp_top.v(481)
    assign n3876 = n3357 ? encrypted_data_buf[1680] : n3868;   // modexp_top.v(481)
    assign n3877 = n3352 ? encrypted_data_buf[1679] : n3869;   // modexp_top.v(481)
    assign n3878 = n3352 ? encrypted_data_buf[1678] : n3870;   // modexp_top.v(481)
    assign n3879 = n3352 ? encrypted_data_buf[1677] : n3871;   // modexp_top.v(481)
    assign n3880 = n3352 ? encrypted_data_buf[1676] : n3872;   // modexp_top.v(481)
    assign n3881 = n3352 ? encrypted_data_buf[1675] : n3873;   // modexp_top.v(481)
    assign n3882 = n3352 ? encrypted_data_buf[1674] : n3874;   // modexp_top.v(481)
    assign n3883 = n3352 ? encrypted_data_buf[1673] : n3875;   // modexp_top.v(481)
    assign n3884 = n3352 ? encrypted_data_buf[1672] : n3876;   // modexp_top.v(481)
    assign n3885 = n3347 ? encrypted_data_buf[1671] : n3877;   // modexp_top.v(481)
    assign n3886 = n3347 ? encrypted_data_buf[1670] : n3878;   // modexp_top.v(481)
    assign n3887 = n3347 ? encrypted_data_buf[1669] : n3879;   // modexp_top.v(481)
    assign n3888 = n3347 ? encrypted_data_buf[1668] : n3880;   // modexp_top.v(481)
    assign n3889 = n3347 ? encrypted_data_buf[1667] : n3881;   // modexp_top.v(481)
    assign n3890 = n3347 ? encrypted_data_buf[1666] : n3882;   // modexp_top.v(481)
    assign n3891 = n3347 ? encrypted_data_buf[1665] : n3883;   // modexp_top.v(481)
    assign n3892 = n3347 ? encrypted_data_buf[1664] : n3884;   // modexp_top.v(481)
    assign n3893 = n3341 ? encrypted_data_buf[1663] : n3885;   // modexp_top.v(481)
    assign n3894 = n3341 ? encrypted_data_buf[1662] : n3886;   // modexp_top.v(481)
    assign n3895 = n3341 ? encrypted_data_buf[1661] : n3887;   // modexp_top.v(481)
    assign n3896 = n3341 ? encrypted_data_buf[1660] : n3888;   // modexp_top.v(481)
    assign n3897 = n3341 ? encrypted_data_buf[1659] : n3889;   // modexp_top.v(481)
    assign n3898 = n3341 ? encrypted_data_buf[1658] : n3890;   // modexp_top.v(481)
    assign n3899 = n3341 ? encrypted_data_buf[1657] : n3891;   // modexp_top.v(481)
    assign n3900 = n3341 ? encrypted_data_buf[1656] : n3892;   // modexp_top.v(481)
    assign n3901 = n3338 ? encrypted_data_buf[1655] : n3893;   // modexp_top.v(481)
    assign n3902 = n3338 ? encrypted_data_buf[1654] : n3894;   // modexp_top.v(481)
    assign n3903 = n3338 ? encrypted_data_buf[1653] : n3895;   // modexp_top.v(481)
    assign n3904 = n3338 ? encrypted_data_buf[1652] : n3896;   // modexp_top.v(481)
    assign n3905 = n3338 ? encrypted_data_buf[1651] : n3897;   // modexp_top.v(481)
    assign n3906 = n3338 ? encrypted_data_buf[1650] : n3898;   // modexp_top.v(481)
    assign n3907 = n3338 ? encrypted_data_buf[1649] : n3899;   // modexp_top.v(481)
    assign n3908 = n3338 ? encrypted_data_buf[1648] : n3900;   // modexp_top.v(481)
    assign n3909 = n3334 ? encrypted_data_buf[1647] : n3901;   // modexp_top.v(481)
    assign n3910 = n3334 ? encrypted_data_buf[1646] : n3902;   // modexp_top.v(481)
    assign n3911 = n3334 ? encrypted_data_buf[1645] : n3903;   // modexp_top.v(481)
    assign n3912 = n3334 ? encrypted_data_buf[1644] : n3904;   // modexp_top.v(481)
    assign n3913 = n3334 ? encrypted_data_buf[1643] : n3905;   // modexp_top.v(481)
    assign n3914 = n3334 ? encrypted_data_buf[1642] : n3906;   // modexp_top.v(481)
    assign n3915 = n3334 ? encrypted_data_buf[1641] : n3907;   // modexp_top.v(481)
    assign n3916 = n3334 ? encrypted_data_buf[1640] : n3908;   // modexp_top.v(481)
    assign n3917 = n3330 ? encrypted_data_buf[1639] : n3909;   // modexp_top.v(481)
    assign n3918 = n3330 ? encrypted_data_buf[1638] : n3910;   // modexp_top.v(481)
    assign n3919 = n3330 ? encrypted_data_buf[1637] : n3911;   // modexp_top.v(481)
    assign n3920 = n3330 ? encrypted_data_buf[1636] : n3912;   // modexp_top.v(481)
    assign n3921 = n3330 ? encrypted_data_buf[1635] : n3913;   // modexp_top.v(481)
    assign n3922 = n3330 ? encrypted_data_buf[1634] : n3914;   // modexp_top.v(481)
    assign n3923 = n3330 ? encrypted_data_buf[1633] : n3915;   // modexp_top.v(481)
    assign n3924 = n3330 ? encrypted_data_buf[1632] : n3916;   // modexp_top.v(481)
    assign n3925 = n3325 ? encrypted_data_buf[1631] : n3917;   // modexp_top.v(481)
    assign n3926 = n3325 ? encrypted_data_buf[1630] : n3918;   // modexp_top.v(481)
    assign n3927 = n3325 ? encrypted_data_buf[1629] : n3919;   // modexp_top.v(481)
    assign n3928 = n3325 ? encrypted_data_buf[1628] : n3920;   // modexp_top.v(481)
    assign n3929 = n3325 ? encrypted_data_buf[1627] : n3921;   // modexp_top.v(481)
    assign n3930 = n3325 ? encrypted_data_buf[1626] : n3922;   // modexp_top.v(481)
    assign n3931 = n3325 ? encrypted_data_buf[1625] : n3923;   // modexp_top.v(481)
    assign n3932 = n3325 ? encrypted_data_buf[1624] : n3924;   // modexp_top.v(481)
    assign n3933 = n3321 ? encrypted_data_buf[1623] : n3925;   // modexp_top.v(481)
    assign n3934 = n3321 ? encrypted_data_buf[1622] : n3926;   // modexp_top.v(481)
    assign n3935 = n3321 ? encrypted_data_buf[1621] : n3927;   // modexp_top.v(481)
    assign n3936 = n3321 ? encrypted_data_buf[1620] : n3928;   // modexp_top.v(481)
    assign n3937 = n3321 ? encrypted_data_buf[1619] : n3929;   // modexp_top.v(481)
    assign n3938 = n3321 ? encrypted_data_buf[1618] : n3930;   // modexp_top.v(481)
    assign n3939 = n3321 ? encrypted_data_buf[1617] : n3931;   // modexp_top.v(481)
    assign n3940 = n3321 ? encrypted_data_buf[1616] : n3932;   // modexp_top.v(481)
    assign n3941 = n3316 ? encrypted_data_buf[1615] : n3933;   // modexp_top.v(481)
    assign n3942 = n3316 ? encrypted_data_buf[1614] : n3934;   // modexp_top.v(481)
    assign n3943 = n3316 ? encrypted_data_buf[1613] : n3935;   // modexp_top.v(481)
    assign n3944 = n3316 ? encrypted_data_buf[1612] : n3936;   // modexp_top.v(481)
    assign n3945 = n3316 ? encrypted_data_buf[1611] : n3937;   // modexp_top.v(481)
    assign n3946 = n3316 ? encrypted_data_buf[1610] : n3938;   // modexp_top.v(481)
    assign n3947 = n3316 ? encrypted_data_buf[1609] : n3939;   // modexp_top.v(481)
    assign n3948 = n3316 ? encrypted_data_buf[1608] : n3940;   // modexp_top.v(481)
    assign n3949 = n3311 ? encrypted_data_buf[1607] : n3941;   // modexp_top.v(481)
    assign n3950 = n3311 ? encrypted_data_buf[1606] : n3942;   // modexp_top.v(481)
    assign n3951 = n3311 ? encrypted_data_buf[1605] : n3943;   // modexp_top.v(481)
    assign n3952 = n3311 ? encrypted_data_buf[1604] : n3944;   // modexp_top.v(481)
    assign n3953 = n3311 ? encrypted_data_buf[1603] : n3945;   // modexp_top.v(481)
    assign n3954 = n3311 ? encrypted_data_buf[1602] : n3946;   // modexp_top.v(481)
    assign n3955 = n3311 ? encrypted_data_buf[1601] : n3947;   // modexp_top.v(481)
    assign n3956 = n3311 ? encrypted_data_buf[1600] : n3948;   // modexp_top.v(481)
    assign n3957 = n3305 ? encrypted_data_buf[1599] : n3949;   // modexp_top.v(481)
    assign n3958 = n3305 ? encrypted_data_buf[1598] : n3950;   // modexp_top.v(481)
    assign n3959 = n3305 ? encrypted_data_buf[1597] : n3951;   // modexp_top.v(481)
    assign n3960 = n3305 ? encrypted_data_buf[1596] : n3952;   // modexp_top.v(481)
    assign n3961 = n3305 ? encrypted_data_buf[1595] : n3953;   // modexp_top.v(481)
    assign n3962 = n3305 ? encrypted_data_buf[1594] : n3954;   // modexp_top.v(481)
    assign n3963 = n3305 ? encrypted_data_buf[1593] : n3955;   // modexp_top.v(481)
    assign n3964 = n3305 ? encrypted_data_buf[1592] : n3956;   // modexp_top.v(481)
    assign n3965 = n3301 ? encrypted_data_buf[1591] : n3957;   // modexp_top.v(481)
    assign n3966 = n3301 ? encrypted_data_buf[1590] : n3958;   // modexp_top.v(481)
    assign n3967 = n3301 ? encrypted_data_buf[1589] : n3959;   // modexp_top.v(481)
    assign n3968 = n3301 ? encrypted_data_buf[1588] : n3960;   // modexp_top.v(481)
    assign n3969 = n3301 ? encrypted_data_buf[1587] : n3961;   // modexp_top.v(481)
    assign n3970 = n3301 ? encrypted_data_buf[1586] : n3962;   // modexp_top.v(481)
    assign n3971 = n3301 ? encrypted_data_buf[1585] : n3963;   // modexp_top.v(481)
    assign n3972 = n3301 ? encrypted_data_buf[1584] : n3964;   // modexp_top.v(481)
    assign n3973 = n3296 ? encrypted_data_buf[1583] : n3965;   // modexp_top.v(481)
    assign n3974 = n3296 ? encrypted_data_buf[1582] : n3966;   // modexp_top.v(481)
    assign n3975 = n3296 ? encrypted_data_buf[1581] : n3967;   // modexp_top.v(481)
    assign n3976 = n3296 ? encrypted_data_buf[1580] : n3968;   // modexp_top.v(481)
    assign n3977 = n3296 ? encrypted_data_buf[1579] : n3969;   // modexp_top.v(481)
    assign n3978 = n3296 ? encrypted_data_buf[1578] : n3970;   // modexp_top.v(481)
    assign n3979 = n3296 ? encrypted_data_buf[1577] : n3971;   // modexp_top.v(481)
    assign n3980 = n3296 ? encrypted_data_buf[1576] : n3972;   // modexp_top.v(481)
    assign n3981 = n3291 ? encrypted_data_buf[1575] : n3973;   // modexp_top.v(481)
    assign n3982 = n3291 ? encrypted_data_buf[1574] : n3974;   // modexp_top.v(481)
    assign n3983 = n3291 ? encrypted_data_buf[1573] : n3975;   // modexp_top.v(481)
    assign n3984 = n3291 ? encrypted_data_buf[1572] : n3976;   // modexp_top.v(481)
    assign n3985 = n3291 ? encrypted_data_buf[1571] : n3977;   // modexp_top.v(481)
    assign n3986 = n3291 ? encrypted_data_buf[1570] : n3978;   // modexp_top.v(481)
    assign n3987 = n3291 ? encrypted_data_buf[1569] : n3979;   // modexp_top.v(481)
    assign n3988 = n3291 ? encrypted_data_buf[1568] : n3980;   // modexp_top.v(481)
    assign n3989 = n3285 ? encrypted_data_buf[1567] : n3981;   // modexp_top.v(481)
    assign n3990 = n3285 ? encrypted_data_buf[1566] : n3982;   // modexp_top.v(481)
    assign n3991 = n3285 ? encrypted_data_buf[1565] : n3983;   // modexp_top.v(481)
    assign n3992 = n3285 ? encrypted_data_buf[1564] : n3984;   // modexp_top.v(481)
    assign n3993 = n3285 ? encrypted_data_buf[1563] : n3985;   // modexp_top.v(481)
    assign n3994 = n3285 ? encrypted_data_buf[1562] : n3986;   // modexp_top.v(481)
    assign n3995 = n3285 ? encrypted_data_buf[1561] : n3987;   // modexp_top.v(481)
    assign n3996 = n3285 ? encrypted_data_buf[1560] : n3988;   // modexp_top.v(481)
    assign n3997 = n3280 ? encrypted_data_buf[1559] : n3989;   // modexp_top.v(481)
    assign n3998 = n3280 ? encrypted_data_buf[1558] : n3990;   // modexp_top.v(481)
    assign n3999 = n3280 ? encrypted_data_buf[1557] : n3991;   // modexp_top.v(481)
    assign n4000 = n3280 ? encrypted_data_buf[1556] : n3992;   // modexp_top.v(481)
    assign n4001 = n3280 ? encrypted_data_buf[1555] : n3993;   // modexp_top.v(481)
    assign n4002 = n3280 ? encrypted_data_buf[1554] : n3994;   // modexp_top.v(481)
    assign n4003 = n3280 ? encrypted_data_buf[1553] : n3995;   // modexp_top.v(481)
    assign n4004 = n3280 ? encrypted_data_buf[1552] : n3996;   // modexp_top.v(481)
    assign n4005 = n3274 ? encrypted_data_buf[1551] : n3997;   // modexp_top.v(481)
    assign n4006 = n3274 ? encrypted_data_buf[1550] : n3998;   // modexp_top.v(481)
    assign n4007 = n3274 ? encrypted_data_buf[1549] : n3999;   // modexp_top.v(481)
    assign n4008 = n3274 ? encrypted_data_buf[1548] : n4000;   // modexp_top.v(481)
    assign n4009 = n3274 ? encrypted_data_buf[1547] : n4001;   // modexp_top.v(481)
    assign n4010 = n3274 ? encrypted_data_buf[1546] : n4002;   // modexp_top.v(481)
    assign n4011 = n3274 ? encrypted_data_buf[1545] : n4003;   // modexp_top.v(481)
    assign n4012 = n3274 ? encrypted_data_buf[1544] : n4004;   // modexp_top.v(481)
    assign n4013 = n3268 ? encrypted_data_buf[1543] : n4005;   // modexp_top.v(481)
    assign n4014 = n3268 ? encrypted_data_buf[1542] : n4006;   // modexp_top.v(481)
    assign n4015 = n3268 ? encrypted_data_buf[1541] : n4007;   // modexp_top.v(481)
    assign n4016 = n3268 ? encrypted_data_buf[1540] : n4008;   // modexp_top.v(481)
    assign n4017 = n3268 ? encrypted_data_buf[1539] : n4009;   // modexp_top.v(481)
    assign n4018 = n3268 ? encrypted_data_buf[1538] : n4010;   // modexp_top.v(481)
    assign n4019 = n3268 ? encrypted_data_buf[1537] : n4011;   // modexp_top.v(481)
    assign n4020 = n3268 ? encrypted_data_buf[1536] : n4012;   // modexp_top.v(481)
    assign n4021 = n3261 ? encrypted_data_buf[1535] : n4013;   // modexp_top.v(481)
    assign n4022 = n3261 ? encrypted_data_buf[1534] : n4014;   // modexp_top.v(481)
    assign n4023 = n3261 ? encrypted_data_buf[1533] : n4015;   // modexp_top.v(481)
    assign n4024 = n3261 ? encrypted_data_buf[1532] : n4016;   // modexp_top.v(481)
    assign n4025 = n3261 ? encrypted_data_buf[1531] : n4017;   // modexp_top.v(481)
    assign n4026 = n3261 ? encrypted_data_buf[1530] : n4018;   // modexp_top.v(481)
    assign n4027 = n3261 ? encrypted_data_buf[1529] : n4019;   // modexp_top.v(481)
    assign n4028 = n3261 ? encrypted_data_buf[1528] : n4020;   // modexp_top.v(481)
    assign n4029 = n3259 ? encrypted_data_buf[1527] : n4021;   // modexp_top.v(481)
    assign n4030 = n3259 ? encrypted_data_buf[1526] : n4022;   // modexp_top.v(481)
    assign n4031 = n3259 ? encrypted_data_buf[1525] : n4023;   // modexp_top.v(481)
    assign n4032 = n3259 ? encrypted_data_buf[1524] : n4024;   // modexp_top.v(481)
    assign n4033 = n3259 ? encrypted_data_buf[1523] : n4025;   // modexp_top.v(481)
    assign n4034 = n3259 ? encrypted_data_buf[1522] : n4026;   // modexp_top.v(481)
    assign n4035 = n3259 ? encrypted_data_buf[1521] : n4027;   // modexp_top.v(481)
    assign n4036 = n3259 ? encrypted_data_buf[1520] : n4028;   // modexp_top.v(481)
    assign n4037 = n3256 ? encrypted_data_buf[1519] : n4029;   // modexp_top.v(481)
    assign n4038 = n3256 ? encrypted_data_buf[1518] : n4030;   // modexp_top.v(481)
    assign n4039 = n3256 ? encrypted_data_buf[1517] : n4031;   // modexp_top.v(481)
    assign n4040 = n3256 ? encrypted_data_buf[1516] : n4032;   // modexp_top.v(481)
    assign n4041 = n3256 ? encrypted_data_buf[1515] : n4033;   // modexp_top.v(481)
    assign n4042 = n3256 ? encrypted_data_buf[1514] : n4034;   // modexp_top.v(481)
    assign n4043 = n3256 ? encrypted_data_buf[1513] : n4035;   // modexp_top.v(481)
    assign n4044 = n3256 ? encrypted_data_buf[1512] : n4036;   // modexp_top.v(481)
    assign n4045 = n3253 ? encrypted_data_buf[1511] : n4037;   // modexp_top.v(481)
    assign n4046 = n3253 ? encrypted_data_buf[1510] : n4038;   // modexp_top.v(481)
    assign n4047 = n3253 ? encrypted_data_buf[1509] : n4039;   // modexp_top.v(481)
    assign n4048 = n3253 ? encrypted_data_buf[1508] : n4040;   // modexp_top.v(481)
    assign n4049 = n3253 ? encrypted_data_buf[1507] : n4041;   // modexp_top.v(481)
    assign n4050 = n3253 ? encrypted_data_buf[1506] : n4042;   // modexp_top.v(481)
    assign n4051 = n3253 ? encrypted_data_buf[1505] : n4043;   // modexp_top.v(481)
    assign n4052 = n3253 ? encrypted_data_buf[1504] : n4044;   // modexp_top.v(481)
    assign n4053 = n3249 ? encrypted_data_buf[1503] : n4045;   // modexp_top.v(481)
    assign n4054 = n3249 ? encrypted_data_buf[1502] : n4046;   // modexp_top.v(481)
    assign n4055 = n3249 ? encrypted_data_buf[1501] : n4047;   // modexp_top.v(481)
    assign n4056 = n3249 ? encrypted_data_buf[1500] : n4048;   // modexp_top.v(481)
    assign n4057 = n3249 ? encrypted_data_buf[1499] : n4049;   // modexp_top.v(481)
    assign n4058 = n3249 ? encrypted_data_buf[1498] : n4050;   // modexp_top.v(481)
    assign n4059 = n3249 ? encrypted_data_buf[1497] : n4051;   // modexp_top.v(481)
    assign n4060 = n3249 ? encrypted_data_buf[1496] : n4052;   // modexp_top.v(481)
    assign n4061 = n3246 ? encrypted_data_buf[1495] : n4053;   // modexp_top.v(481)
    assign n4062 = n3246 ? encrypted_data_buf[1494] : n4054;   // modexp_top.v(481)
    assign n4063 = n3246 ? encrypted_data_buf[1493] : n4055;   // modexp_top.v(481)
    assign n4064 = n3246 ? encrypted_data_buf[1492] : n4056;   // modexp_top.v(481)
    assign n4065 = n3246 ? encrypted_data_buf[1491] : n4057;   // modexp_top.v(481)
    assign n4066 = n3246 ? encrypted_data_buf[1490] : n4058;   // modexp_top.v(481)
    assign n4067 = n3246 ? encrypted_data_buf[1489] : n4059;   // modexp_top.v(481)
    assign n4068 = n3246 ? encrypted_data_buf[1488] : n4060;   // modexp_top.v(481)
    assign n4069 = n3242 ? encrypted_data_buf[1487] : n4061;   // modexp_top.v(481)
    assign n4070 = n3242 ? encrypted_data_buf[1486] : n4062;   // modexp_top.v(481)
    assign n4071 = n3242 ? encrypted_data_buf[1485] : n4063;   // modexp_top.v(481)
    assign n4072 = n3242 ? encrypted_data_buf[1484] : n4064;   // modexp_top.v(481)
    assign n4073 = n3242 ? encrypted_data_buf[1483] : n4065;   // modexp_top.v(481)
    assign n4074 = n3242 ? encrypted_data_buf[1482] : n4066;   // modexp_top.v(481)
    assign n4075 = n3242 ? encrypted_data_buf[1481] : n4067;   // modexp_top.v(481)
    assign n4076 = n3242 ? encrypted_data_buf[1480] : n4068;   // modexp_top.v(481)
    assign n4077 = n3238 ? encrypted_data_buf[1479] : n4069;   // modexp_top.v(481)
    assign n4078 = n3238 ? encrypted_data_buf[1478] : n4070;   // modexp_top.v(481)
    assign n4079 = n3238 ? encrypted_data_buf[1477] : n4071;   // modexp_top.v(481)
    assign n4080 = n3238 ? encrypted_data_buf[1476] : n4072;   // modexp_top.v(481)
    assign n4081 = n3238 ? encrypted_data_buf[1475] : n4073;   // modexp_top.v(481)
    assign n4082 = n3238 ? encrypted_data_buf[1474] : n4074;   // modexp_top.v(481)
    assign n4083 = n3238 ? encrypted_data_buf[1473] : n4075;   // modexp_top.v(481)
    assign n4084 = n3238 ? encrypted_data_buf[1472] : n4076;   // modexp_top.v(481)
    assign n4085 = n3233 ? encrypted_data_buf[1471] : n4077;   // modexp_top.v(481)
    assign n4086 = n3233 ? encrypted_data_buf[1470] : n4078;   // modexp_top.v(481)
    assign n4087 = n3233 ? encrypted_data_buf[1469] : n4079;   // modexp_top.v(481)
    assign n4088 = n3233 ? encrypted_data_buf[1468] : n4080;   // modexp_top.v(481)
    assign n4089 = n3233 ? encrypted_data_buf[1467] : n4081;   // modexp_top.v(481)
    assign n4090 = n3233 ? encrypted_data_buf[1466] : n4082;   // modexp_top.v(481)
    assign n4091 = n3233 ? encrypted_data_buf[1465] : n4083;   // modexp_top.v(481)
    assign n4092 = n3233 ? encrypted_data_buf[1464] : n4084;   // modexp_top.v(481)
    assign n4093 = n3230 ? encrypted_data_buf[1463] : n4085;   // modexp_top.v(481)
    assign n4094 = n3230 ? encrypted_data_buf[1462] : n4086;   // modexp_top.v(481)
    assign n4095 = n3230 ? encrypted_data_buf[1461] : n4087;   // modexp_top.v(481)
    assign n4096 = n3230 ? encrypted_data_buf[1460] : n4088;   // modexp_top.v(481)
    assign n4097 = n3230 ? encrypted_data_buf[1459] : n4089;   // modexp_top.v(481)
    assign n4098 = n3230 ? encrypted_data_buf[1458] : n4090;   // modexp_top.v(481)
    assign n4099 = n3230 ? encrypted_data_buf[1457] : n4091;   // modexp_top.v(481)
    assign n4100 = n3230 ? encrypted_data_buf[1456] : n4092;   // modexp_top.v(481)
    assign n4101 = n3226 ? encrypted_data_buf[1455] : n4093;   // modexp_top.v(481)
    assign n4102 = n3226 ? encrypted_data_buf[1454] : n4094;   // modexp_top.v(481)
    assign n4103 = n3226 ? encrypted_data_buf[1453] : n4095;   // modexp_top.v(481)
    assign n4104 = n3226 ? encrypted_data_buf[1452] : n4096;   // modexp_top.v(481)
    assign n4105 = n3226 ? encrypted_data_buf[1451] : n4097;   // modexp_top.v(481)
    assign n4106 = n3226 ? encrypted_data_buf[1450] : n4098;   // modexp_top.v(481)
    assign n4107 = n3226 ? encrypted_data_buf[1449] : n4099;   // modexp_top.v(481)
    assign n4108 = n3226 ? encrypted_data_buf[1448] : n4100;   // modexp_top.v(481)
    assign n4109 = n3222 ? encrypted_data_buf[1447] : n4101;   // modexp_top.v(481)
    assign n4110 = n3222 ? encrypted_data_buf[1446] : n4102;   // modexp_top.v(481)
    assign n4111 = n3222 ? encrypted_data_buf[1445] : n4103;   // modexp_top.v(481)
    assign n4112 = n3222 ? encrypted_data_buf[1444] : n4104;   // modexp_top.v(481)
    assign n4113 = n3222 ? encrypted_data_buf[1443] : n4105;   // modexp_top.v(481)
    assign n4114 = n3222 ? encrypted_data_buf[1442] : n4106;   // modexp_top.v(481)
    assign n4115 = n3222 ? encrypted_data_buf[1441] : n4107;   // modexp_top.v(481)
    assign n4116 = n3222 ? encrypted_data_buf[1440] : n4108;   // modexp_top.v(481)
    assign n4117 = n3217 ? encrypted_data_buf[1439] : n4109;   // modexp_top.v(481)
    assign n4118 = n3217 ? encrypted_data_buf[1438] : n4110;   // modexp_top.v(481)
    assign n4119 = n3217 ? encrypted_data_buf[1437] : n4111;   // modexp_top.v(481)
    assign n4120 = n3217 ? encrypted_data_buf[1436] : n4112;   // modexp_top.v(481)
    assign n4121 = n3217 ? encrypted_data_buf[1435] : n4113;   // modexp_top.v(481)
    assign n4122 = n3217 ? encrypted_data_buf[1434] : n4114;   // modexp_top.v(481)
    assign n4123 = n3217 ? encrypted_data_buf[1433] : n4115;   // modexp_top.v(481)
    assign n4124 = n3217 ? encrypted_data_buf[1432] : n4116;   // modexp_top.v(481)
    assign n4125 = n3213 ? encrypted_data_buf[1431] : n4117;   // modexp_top.v(481)
    assign n4126 = n3213 ? encrypted_data_buf[1430] : n4118;   // modexp_top.v(481)
    assign n4127 = n3213 ? encrypted_data_buf[1429] : n4119;   // modexp_top.v(481)
    assign n4128 = n3213 ? encrypted_data_buf[1428] : n4120;   // modexp_top.v(481)
    assign n4129 = n3213 ? encrypted_data_buf[1427] : n4121;   // modexp_top.v(481)
    assign n4130 = n3213 ? encrypted_data_buf[1426] : n4122;   // modexp_top.v(481)
    assign n4131 = n3213 ? encrypted_data_buf[1425] : n4123;   // modexp_top.v(481)
    assign n4132 = n3213 ? encrypted_data_buf[1424] : n4124;   // modexp_top.v(481)
    assign n4133 = n3208 ? encrypted_data_buf[1423] : n4125;   // modexp_top.v(481)
    assign n4134 = n3208 ? encrypted_data_buf[1422] : n4126;   // modexp_top.v(481)
    assign n4135 = n3208 ? encrypted_data_buf[1421] : n4127;   // modexp_top.v(481)
    assign n4136 = n3208 ? encrypted_data_buf[1420] : n4128;   // modexp_top.v(481)
    assign n4137 = n3208 ? encrypted_data_buf[1419] : n4129;   // modexp_top.v(481)
    assign n4138 = n3208 ? encrypted_data_buf[1418] : n4130;   // modexp_top.v(481)
    assign n4139 = n3208 ? encrypted_data_buf[1417] : n4131;   // modexp_top.v(481)
    assign n4140 = n3208 ? encrypted_data_buf[1416] : n4132;   // modexp_top.v(481)
    assign n4141 = n3203 ? encrypted_data_buf[1415] : n4133;   // modexp_top.v(481)
    assign n4142 = n3203 ? encrypted_data_buf[1414] : n4134;   // modexp_top.v(481)
    assign n4143 = n3203 ? encrypted_data_buf[1413] : n4135;   // modexp_top.v(481)
    assign n4144 = n3203 ? encrypted_data_buf[1412] : n4136;   // modexp_top.v(481)
    assign n4145 = n3203 ? encrypted_data_buf[1411] : n4137;   // modexp_top.v(481)
    assign n4146 = n3203 ? encrypted_data_buf[1410] : n4138;   // modexp_top.v(481)
    assign n4147 = n3203 ? encrypted_data_buf[1409] : n4139;   // modexp_top.v(481)
    assign n4148 = n3203 ? encrypted_data_buf[1408] : n4140;   // modexp_top.v(481)
    assign n4149 = n3197 ? encrypted_data_buf[1407] : n4141;   // modexp_top.v(481)
    assign n4150 = n3197 ? encrypted_data_buf[1406] : n4142;   // modexp_top.v(481)
    assign n4151 = n3197 ? encrypted_data_buf[1405] : n4143;   // modexp_top.v(481)
    assign n4152 = n3197 ? encrypted_data_buf[1404] : n4144;   // modexp_top.v(481)
    assign n4153 = n3197 ? encrypted_data_buf[1403] : n4145;   // modexp_top.v(481)
    assign n4154 = n3197 ? encrypted_data_buf[1402] : n4146;   // modexp_top.v(481)
    assign n4155 = n3197 ? encrypted_data_buf[1401] : n4147;   // modexp_top.v(481)
    assign n4156 = n3197 ? encrypted_data_buf[1400] : n4148;   // modexp_top.v(481)
    assign n4157 = n3194 ? encrypted_data_buf[1399] : n4149;   // modexp_top.v(481)
    assign n4158 = n3194 ? encrypted_data_buf[1398] : n4150;   // modexp_top.v(481)
    assign n4159 = n3194 ? encrypted_data_buf[1397] : n4151;   // modexp_top.v(481)
    assign n4160 = n3194 ? encrypted_data_buf[1396] : n4152;   // modexp_top.v(481)
    assign n4161 = n3194 ? encrypted_data_buf[1395] : n4153;   // modexp_top.v(481)
    assign n4162 = n3194 ? encrypted_data_buf[1394] : n4154;   // modexp_top.v(481)
    assign n4163 = n3194 ? encrypted_data_buf[1393] : n4155;   // modexp_top.v(481)
    assign n4164 = n3194 ? encrypted_data_buf[1392] : n4156;   // modexp_top.v(481)
    assign n4165 = n3190 ? encrypted_data_buf[1391] : n4157;   // modexp_top.v(481)
    assign n4166 = n3190 ? encrypted_data_buf[1390] : n4158;   // modexp_top.v(481)
    assign n4167 = n3190 ? encrypted_data_buf[1389] : n4159;   // modexp_top.v(481)
    assign n4168 = n3190 ? encrypted_data_buf[1388] : n4160;   // modexp_top.v(481)
    assign n4169 = n3190 ? encrypted_data_buf[1387] : n4161;   // modexp_top.v(481)
    assign n4170 = n3190 ? encrypted_data_buf[1386] : n4162;   // modexp_top.v(481)
    assign n4171 = n3190 ? encrypted_data_buf[1385] : n4163;   // modexp_top.v(481)
    assign n4172 = n3190 ? encrypted_data_buf[1384] : n4164;   // modexp_top.v(481)
    assign n4173 = n3186 ? encrypted_data_buf[1383] : n4165;   // modexp_top.v(481)
    assign n4174 = n3186 ? encrypted_data_buf[1382] : n4166;   // modexp_top.v(481)
    assign n4175 = n3186 ? encrypted_data_buf[1381] : n4167;   // modexp_top.v(481)
    assign n4176 = n3186 ? encrypted_data_buf[1380] : n4168;   // modexp_top.v(481)
    assign n4177 = n3186 ? encrypted_data_buf[1379] : n4169;   // modexp_top.v(481)
    assign n4178 = n3186 ? encrypted_data_buf[1378] : n4170;   // modexp_top.v(481)
    assign n4179 = n3186 ? encrypted_data_buf[1377] : n4171;   // modexp_top.v(481)
    assign n4180 = n3186 ? encrypted_data_buf[1376] : n4172;   // modexp_top.v(481)
    assign n4181 = n3181 ? encrypted_data_buf[1375] : n4173;   // modexp_top.v(481)
    assign n4182 = n3181 ? encrypted_data_buf[1374] : n4174;   // modexp_top.v(481)
    assign n4183 = n3181 ? encrypted_data_buf[1373] : n4175;   // modexp_top.v(481)
    assign n4184 = n3181 ? encrypted_data_buf[1372] : n4176;   // modexp_top.v(481)
    assign n4185 = n3181 ? encrypted_data_buf[1371] : n4177;   // modexp_top.v(481)
    assign n4186 = n3181 ? encrypted_data_buf[1370] : n4178;   // modexp_top.v(481)
    assign n4187 = n3181 ? encrypted_data_buf[1369] : n4179;   // modexp_top.v(481)
    assign n4188 = n3181 ? encrypted_data_buf[1368] : n4180;   // modexp_top.v(481)
    assign n4189 = n3177 ? encrypted_data_buf[1367] : n4181;   // modexp_top.v(481)
    assign n4190 = n3177 ? encrypted_data_buf[1366] : n4182;   // modexp_top.v(481)
    assign n4191 = n3177 ? encrypted_data_buf[1365] : n4183;   // modexp_top.v(481)
    assign n4192 = n3177 ? encrypted_data_buf[1364] : n4184;   // modexp_top.v(481)
    assign n4193 = n3177 ? encrypted_data_buf[1363] : n4185;   // modexp_top.v(481)
    assign n4194 = n3177 ? encrypted_data_buf[1362] : n4186;   // modexp_top.v(481)
    assign n4195 = n3177 ? encrypted_data_buf[1361] : n4187;   // modexp_top.v(481)
    assign n4196 = n3177 ? encrypted_data_buf[1360] : n4188;   // modexp_top.v(481)
    assign n4197 = n3172 ? encrypted_data_buf[1359] : n4189;   // modexp_top.v(481)
    assign n4198 = n3172 ? encrypted_data_buf[1358] : n4190;   // modexp_top.v(481)
    assign n4199 = n3172 ? encrypted_data_buf[1357] : n4191;   // modexp_top.v(481)
    assign n4200 = n3172 ? encrypted_data_buf[1356] : n4192;   // modexp_top.v(481)
    assign n4201 = n3172 ? encrypted_data_buf[1355] : n4193;   // modexp_top.v(481)
    assign n4202 = n3172 ? encrypted_data_buf[1354] : n4194;   // modexp_top.v(481)
    assign n4203 = n3172 ? encrypted_data_buf[1353] : n4195;   // modexp_top.v(481)
    assign n4204 = n3172 ? encrypted_data_buf[1352] : n4196;   // modexp_top.v(481)
    assign n4205 = n3167 ? encrypted_data_buf[1351] : n4197;   // modexp_top.v(481)
    assign n4206 = n3167 ? encrypted_data_buf[1350] : n4198;   // modexp_top.v(481)
    assign n4207 = n3167 ? encrypted_data_buf[1349] : n4199;   // modexp_top.v(481)
    assign n4208 = n3167 ? encrypted_data_buf[1348] : n4200;   // modexp_top.v(481)
    assign n4209 = n3167 ? encrypted_data_buf[1347] : n4201;   // modexp_top.v(481)
    assign n4210 = n3167 ? encrypted_data_buf[1346] : n4202;   // modexp_top.v(481)
    assign n4211 = n3167 ? encrypted_data_buf[1345] : n4203;   // modexp_top.v(481)
    assign n4212 = n3167 ? encrypted_data_buf[1344] : n4204;   // modexp_top.v(481)
    assign n4213 = n3161 ? encrypted_data_buf[1343] : n4205;   // modexp_top.v(481)
    assign n4214 = n3161 ? encrypted_data_buf[1342] : n4206;   // modexp_top.v(481)
    assign n4215 = n3161 ? encrypted_data_buf[1341] : n4207;   // modexp_top.v(481)
    assign n4216 = n3161 ? encrypted_data_buf[1340] : n4208;   // modexp_top.v(481)
    assign n4217 = n3161 ? encrypted_data_buf[1339] : n4209;   // modexp_top.v(481)
    assign n4218 = n3161 ? encrypted_data_buf[1338] : n4210;   // modexp_top.v(481)
    assign n4219 = n3161 ? encrypted_data_buf[1337] : n4211;   // modexp_top.v(481)
    assign n4220 = n3161 ? encrypted_data_buf[1336] : n4212;   // modexp_top.v(481)
    assign n4221 = n3157 ? encrypted_data_buf[1335] : n4213;   // modexp_top.v(481)
    assign n4222 = n3157 ? encrypted_data_buf[1334] : n4214;   // modexp_top.v(481)
    assign n4223 = n3157 ? encrypted_data_buf[1333] : n4215;   // modexp_top.v(481)
    assign n4224 = n3157 ? encrypted_data_buf[1332] : n4216;   // modexp_top.v(481)
    assign n4225 = n3157 ? encrypted_data_buf[1331] : n4217;   // modexp_top.v(481)
    assign n4226 = n3157 ? encrypted_data_buf[1330] : n4218;   // modexp_top.v(481)
    assign n4227 = n3157 ? encrypted_data_buf[1329] : n4219;   // modexp_top.v(481)
    assign n4228 = n3157 ? encrypted_data_buf[1328] : n4220;   // modexp_top.v(481)
    assign n4229 = n3152 ? encrypted_data_buf[1327] : n4221;   // modexp_top.v(481)
    assign n4230 = n3152 ? encrypted_data_buf[1326] : n4222;   // modexp_top.v(481)
    assign n4231 = n3152 ? encrypted_data_buf[1325] : n4223;   // modexp_top.v(481)
    assign n4232 = n3152 ? encrypted_data_buf[1324] : n4224;   // modexp_top.v(481)
    assign n4233 = n3152 ? encrypted_data_buf[1323] : n4225;   // modexp_top.v(481)
    assign n4234 = n3152 ? encrypted_data_buf[1322] : n4226;   // modexp_top.v(481)
    assign n4235 = n3152 ? encrypted_data_buf[1321] : n4227;   // modexp_top.v(481)
    assign n4236 = n3152 ? encrypted_data_buf[1320] : n4228;   // modexp_top.v(481)
    assign n4237 = n3147 ? encrypted_data_buf[1319] : n4229;   // modexp_top.v(481)
    assign n4238 = n3147 ? encrypted_data_buf[1318] : n4230;   // modexp_top.v(481)
    assign n4239 = n3147 ? encrypted_data_buf[1317] : n4231;   // modexp_top.v(481)
    assign n4240 = n3147 ? encrypted_data_buf[1316] : n4232;   // modexp_top.v(481)
    assign n4241 = n3147 ? encrypted_data_buf[1315] : n4233;   // modexp_top.v(481)
    assign n4242 = n3147 ? encrypted_data_buf[1314] : n4234;   // modexp_top.v(481)
    assign n4243 = n3147 ? encrypted_data_buf[1313] : n4235;   // modexp_top.v(481)
    assign n4244 = n3147 ? encrypted_data_buf[1312] : n4236;   // modexp_top.v(481)
    assign n4245 = n3141 ? encrypted_data_buf[1311] : n4237;   // modexp_top.v(481)
    assign n4246 = n3141 ? encrypted_data_buf[1310] : n4238;   // modexp_top.v(481)
    assign n4247 = n3141 ? encrypted_data_buf[1309] : n4239;   // modexp_top.v(481)
    assign n4248 = n3141 ? encrypted_data_buf[1308] : n4240;   // modexp_top.v(481)
    assign n4249 = n3141 ? encrypted_data_buf[1307] : n4241;   // modexp_top.v(481)
    assign n4250 = n3141 ? encrypted_data_buf[1306] : n4242;   // modexp_top.v(481)
    assign n4251 = n3141 ? encrypted_data_buf[1305] : n4243;   // modexp_top.v(481)
    assign n4252 = n3141 ? encrypted_data_buf[1304] : n4244;   // modexp_top.v(481)
    assign n4253 = n3136 ? encrypted_data_buf[1303] : n4245;   // modexp_top.v(481)
    assign n4254 = n3136 ? encrypted_data_buf[1302] : n4246;   // modexp_top.v(481)
    assign n4255 = n3136 ? encrypted_data_buf[1301] : n4247;   // modexp_top.v(481)
    assign n4256 = n3136 ? encrypted_data_buf[1300] : n4248;   // modexp_top.v(481)
    assign n4257 = n3136 ? encrypted_data_buf[1299] : n4249;   // modexp_top.v(481)
    assign n4258 = n3136 ? encrypted_data_buf[1298] : n4250;   // modexp_top.v(481)
    assign n4259 = n3136 ? encrypted_data_buf[1297] : n4251;   // modexp_top.v(481)
    assign n4260 = n3136 ? encrypted_data_buf[1296] : n4252;   // modexp_top.v(481)
    assign n4261 = n3130 ? encrypted_data_buf[1295] : n4253;   // modexp_top.v(481)
    assign n4262 = n3130 ? encrypted_data_buf[1294] : n4254;   // modexp_top.v(481)
    assign n4263 = n3130 ? encrypted_data_buf[1293] : n4255;   // modexp_top.v(481)
    assign n4264 = n3130 ? encrypted_data_buf[1292] : n4256;   // modexp_top.v(481)
    assign n4265 = n3130 ? encrypted_data_buf[1291] : n4257;   // modexp_top.v(481)
    assign n4266 = n3130 ? encrypted_data_buf[1290] : n4258;   // modexp_top.v(481)
    assign n4267 = n3130 ? encrypted_data_buf[1289] : n4259;   // modexp_top.v(481)
    assign n4268 = n3130 ? encrypted_data_buf[1288] : n4260;   // modexp_top.v(481)
    assign n4269 = n3124 ? encrypted_data_buf[1287] : n4261;   // modexp_top.v(481)
    assign n4270 = n3124 ? encrypted_data_buf[1286] : n4262;   // modexp_top.v(481)
    assign n4271 = n3124 ? encrypted_data_buf[1285] : n4263;   // modexp_top.v(481)
    assign n4272 = n3124 ? encrypted_data_buf[1284] : n4264;   // modexp_top.v(481)
    assign n4273 = n3124 ? encrypted_data_buf[1283] : n4265;   // modexp_top.v(481)
    assign n4274 = n3124 ? encrypted_data_buf[1282] : n4266;   // modexp_top.v(481)
    assign n4275 = n3124 ? encrypted_data_buf[1281] : n4267;   // modexp_top.v(481)
    assign n4276 = n3124 ? encrypted_data_buf[1280] : n4268;   // modexp_top.v(481)
    assign n4277 = n3117 ? encrypted_data_buf[1279] : n4269;   // modexp_top.v(481)
    assign n4278 = n3117 ? encrypted_data_buf[1278] : n4270;   // modexp_top.v(481)
    assign n4279 = n3117 ? encrypted_data_buf[1277] : n4271;   // modexp_top.v(481)
    assign n4280 = n3117 ? encrypted_data_buf[1276] : n4272;   // modexp_top.v(481)
    assign n4281 = n3117 ? encrypted_data_buf[1275] : n4273;   // modexp_top.v(481)
    assign n4282 = n3117 ? encrypted_data_buf[1274] : n4274;   // modexp_top.v(481)
    assign n4283 = n3117 ? encrypted_data_buf[1273] : n4275;   // modexp_top.v(481)
    assign n4284 = n3117 ? encrypted_data_buf[1272] : n4276;   // modexp_top.v(481)
    assign n4285 = n3114 ? encrypted_data_buf[1271] : n4277;   // modexp_top.v(481)
    assign n4286 = n3114 ? encrypted_data_buf[1270] : n4278;   // modexp_top.v(481)
    assign n4287 = n3114 ? encrypted_data_buf[1269] : n4279;   // modexp_top.v(481)
    assign n4288 = n3114 ? encrypted_data_buf[1268] : n4280;   // modexp_top.v(481)
    assign n4289 = n3114 ? encrypted_data_buf[1267] : n4281;   // modexp_top.v(481)
    assign n4290 = n3114 ? encrypted_data_buf[1266] : n4282;   // modexp_top.v(481)
    assign n4291 = n3114 ? encrypted_data_buf[1265] : n4283;   // modexp_top.v(481)
    assign n4292 = n3114 ? encrypted_data_buf[1264] : n4284;   // modexp_top.v(481)
    assign n4293 = n3110 ? encrypted_data_buf[1263] : n4285;   // modexp_top.v(481)
    assign n4294 = n3110 ? encrypted_data_buf[1262] : n4286;   // modexp_top.v(481)
    assign n4295 = n3110 ? encrypted_data_buf[1261] : n4287;   // modexp_top.v(481)
    assign n4296 = n3110 ? encrypted_data_buf[1260] : n4288;   // modexp_top.v(481)
    assign n4297 = n3110 ? encrypted_data_buf[1259] : n4289;   // modexp_top.v(481)
    assign n4298 = n3110 ? encrypted_data_buf[1258] : n4290;   // modexp_top.v(481)
    assign n4299 = n3110 ? encrypted_data_buf[1257] : n4291;   // modexp_top.v(481)
    assign n4300 = n3110 ? encrypted_data_buf[1256] : n4292;   // modexp_top.v(481)
    assign n4301 = n3106 ? encrypted_data_buf[1255] : n4293;   // modexp_top.v(481)
    assign n4302 = n3106 ? encrypted_data_buf[1254] : n4294;   // modexp_top.v(481)
    assign n4303 = n3106 ? encrypted_data_buf[1253] : n4295;   // modexp_top.v(481)
    assign n4304 = n3106 ? encrypted_data_buf[1252] : n4296;   // modexp_top.v(481)
    assign n4305 = n3106 ? encrypted_data_buf[1251] : n4297;   // modexp_top.v(481)
    assign n4306 = n3106 ? encrypted_data_buf[1250] : n4298;   // modexp_top.v(481)
    assign n4307 = n3106 ? encrypted_data_buf[1249] : n4299;   // modexp_top.v(481)
    assign n4308 = n3106 ? encrypted_data_buf[1248] : n4300;   // modexp_top.v(481)
    assign n4309 = n3101 ? encrypted_data_buf[1247] : n4301;   // modexp_top.v(481)
    assign n4310 = n3101 ? encrypted_data_buf[1246] : n4302;   // modexp_top.v(481)
    assign n4311 = n3101 ? encrypted_data_buf[1245] : n4303;   // modexp_top.v(481)
    assign n4312 = n3101 ? encrypted_data_buf[1244] : n4304;   // modexp_top.v(481)
    assign n4313 = n3101 ? encrypted_data_buf[1243] : n4305;   // modexp_top.v(481)
    assign n4314 = n3101 ? encrypted_data_buf[1242] : n4306;   // modexp_top.v(481)
    assign n4315 = n3101 ? encrypted_data_buf[1241] : n4307;   // modexp_top.v(481)
    assign n4316 = n3101 ? encrypted_data_buf[1240] : n4308;   // modexp_top.v(481)
    assign n4317 = n3097 ? encrypted_data_buf[1239] : n4309;   // modexp_top.v(481)
    assign n4318 = n3097 ? encrypted_data_buf[1238] : n4310;   // modexp_top.v(481)
    assign n4319 = n3097 ? encrypted_data_buf[1237] : n4311;   // modexp_top.v(481)
    assign n4320 = n3097 ? encrypted_data_buf[1236] : n4312;   // modexp_top.v(481)
    assign n4321 = n3097 ? encrypted_data_buf[1235] : n4313;   // modexp_top.v(481)
    assign n4322 = n3097 ? encrypted_data_buf[1234] : n4314;   // modexp_top.v(481)
    assign n4323 = n3097 ? encrypted_data_buf[1233] : n4315;   // modexp_top.v(481)
    assign n4324 = n3097 ? encrypted_data_buf[1232] : n4316;   // modexp_top.v(481)
    assign n4325 = n3092 ? encrypted_data_buf[1231] : n4317;   // modexp_top.v(481)
    assign n4326 = n3092 ? encrypted_data_buf[1230] : n4318;   // modexp_top.v(481)
    assign n4327 = n3092 ? encrypted_data_buf[1229] : n4319;   // modexp_top.v(481)
    assign n4328 = n3092 ? encrypted_data_buf[1228] : n4320;   // modexp_top.v(481)
    assign n4329 = n3092 ? encrypted_data_buf[1227] : n4321;   // modexp_top.v(481)
    assign n4330 = n3092 ? encrypted_data_buf[1226] : n4322;   // modexp_top.v(481)
    assign n4331 = n3092 ? encrypted_data_buf[1225] : n4323;   // modexp_top.v(481)
    assign n4332 = n3092 ? encrypted_data_buf[1224] : n4324;   // modexp_top.v(481)
    assign n4333 = n3087 ? encrypted_data_buf[1223] : n4325;   // modexp_top.v(481)
    assign n4334 = n3087 ? encrypted_data_buf[1222] : n4326;   // modexp_top.v(481)
    assign n4335 = n3087 ? encrypted_data_buf[1221] : n4327;   // modexp_top.v(481)
    assign n4336 = n3087 ? encrypted_data_buf[1220] : n4328;   // modexp_top.v(481)
    assign n4337 = n3087 ? encrypted_data_buf[1219] : n4329;   // modexp_top.v(481)
    assign n4338 = n3087 ? encrypted_data_buf[1218] : n4330;   // modexp_top.v(481)
    assign n4339 = n3087 ? encrypted_data_buf[1217] : n4331;   // modexp_top.v(481)
    assign n4340 = n3087 ? encrypted_data_buf[1216] : n4332;   // modexp_top.v(481)
    assign n4341 = n3081 ? encrypted_data_buf[1215] : n4333;   // modexp_top.v(481)
    assign n4342 = n3081 ? encrypted_data_buf[1214] : n4334;   // modexp_top.v(481)
    assign n4343 = n3081 ? encrypted_data_buf[1213] : n4335;   // modexp_top.v(481)
    assign n4344 = n3081 ? encrypted_data_buf[1212] : n4336;   // modexp_top.v(481)
    assign n4345 = n3081 ? encrypted_data_buf[1211] : n4337;   // modexp_top.v(481)
    assign n4346 = n3081 ? encrypted_data_buf[1210] : n4338;   // modexp_top.v(481)
    assign n4347 = n3081 ? encrypted_data_buf[1209] : n4339;   // modexp_top.v(481)
    assign n4348 = n3081 ? encrypted_data_buf[1208] : n4340;   // modexp_top.v(481)
    assign n4349 = n3077 ? encrypted_data_buf[1207] : n4341;   // modexp_top.v(481)
    assign n4350 = n3077 ? encrypted_data_buf[1206] : n4342;   // modexp_top.v(481)
    assign n4351 = n3077 ? encrypted_data_buf[1205] : n4343;   // modexp_top.v(481)
    assign n4352 = n3077 ? encrypted_data_buf[1204] : n4344;   // modexp_top.v(481)
    assign n4353 = n3077 ? encrypted_data_buf[1203] : n4345;   // modexp_top.v(481)
    assign n4354 = n3077 ? encrypted_data_buf[1202] : n4346;   // modexp_top.v(481)
    assign n4355 = n3077 ? encrypted_data_buf[1201] : n4347;   // modexp_top.v(481)
    assign n4356 = n3077 ? encrypted_data_buf[1200] : n4348;   // modexp_top.v(481)
    assign n4357 = n3072 ? encrypted_data_buf[1199] : n4349;   // modexp_top.v(481)
    assign n4358 = n3072 ? encrypted_data_buf[1198] : n4350;   // modexp_top.v(481)
    assign n4359 = n3072 ? encrypted_data_buf[1197] : n4351;   // modexp_top.v(481)
    assign n4360 = n3072 ? encrypted_data_buf[1196] : n4352;   // modexp_top.v(481)
    assign n4361 = n3072 ? encrypted_data_buf[1195] : n4353;   // modexp_top.v(481)
    assign n4362 = n3072 ? encrypted_data_buf[1194] : n4354;   // modexp_top.v(481)
    assign n4363 = n3072 ? encrypted_data_buf[1193] : n4355;   // modexp_top.v(481)
    assign n4364 = n3072 ? encrypted_data_buf[1192] : n4356;   // modexp_top.v(481)
    assign n4365 = n3067 ? encrypted_data_buf[1191] : n4357;   // modexp_top.v(481)
    assign n4366 = n3067 ? encrypted_data_buf[1190] : n4358;   // modexp_top.v(481)
    assign n4367 = n3067 ? encrypted_data_buf[1189] : n4359;   // modexp_top.v(481)
    assign n4368 = n3067 ? encrypted_data_buf[1188] : n4360;   // modexp_top.v(481)
    assign n4369 = n3067 ? encrypted_data_buf[1187] : n4361;   // modexp_top.v(481)
    assign n4370 = n3067 ? encrypted_data_buf[1186] : n4362;   // modexp_top.v(481)
    assign n4371 = n3067 ? encrypted_data_buf[1185] : n4363;   // modexp_top.v(481)
    assign n4372 = n3067 ? encrypted_data_buf[1184] : n4364;   // modexp_top.v(481)
    assign n4373 = n3061 ? encrypted_data_buf[1183] : n4365;   // modexp_top.v(481)
    assign n4374 = n3061 ? encrypted_data_buf[1182] : n4366;   // modexp_top.v(481)
    assign n4375 = n3061 ? encrypted_data_buf[1181] : n4367;   // modexp_top.v(481)
    assign n4376 = n3061 ? encrypted_data_buf[1180] : n4368;   // modexp_top.v(481)
    assign n4377 = n3061 ? encrypted_data_buf[1179] : n4369;   // modexp_top.v(481)
    assign n4378 = n3061 ? encrypted_data_buf[1178] : n4370;   // modexp_top.v(481)
    assign n4379 = n3061 ? encrypted_data_buf[1177] : n4371;   // modexp_top.v(481)
    assign n4380 = n3061 ? encrypted_data_buf[1176] : n4372;   // modexp_top.v(481)
    assign n4381 = n3056 ? encrypted_data_buf[1175] : n4373;   // modexp_top.v(481)
    assign n4382 = n3056 ? encrypted_data_buf[1174] : n4374;   // modexp_top.v(481)
    assign n4383 = n3056 ? encrypted_data_buf[1173] : n4375;   // modexp_top.v(481)
    assign n4384 = n3056 ? encrypted_data_buf[1172] : n4376;   // modexp_top.v(481)
    assign n4385 = n3056 ? encrypted_data_buf[1171] : n4377;   // modexp_top.v(481)
    assign n4386 = n3056 ? encrypted_data_buf[1170] : n4378;   // modexp_top.v(481)
    assign n4387 = n3056 ? encrypted_data_buf[1169] : n4379;   // modexp_top.v(481)
    assign n4388 = n3056 ? encrypted_data_buf[1168] : n4380;   // modexp_top.v(481)
    assign n4389 = n3050 ? encrypted_data_buf[1167] : n4381;   // modexp_top.v(481)
    assign n4390 = n3050 ? encrypted_data_buf[1166] : n4382;   // modexp_top.v(481)
    assign n4391 = n3050 ? encrypted_data_buf[1165] : n4383;   // modexp_top.v(481)
    assign n4392 = n3050 ? encrypted_data_buf[1164] : n4384;   // modexp_top.v(481)
    assign n4393 = n3050 ? encrypted_data_buf[1163] : n4385;   // modexp_top.v(481)
    assign n4394 = n3050 ? encrypted_data_buf[1162] : n4386;   // modexp_top.v(481)
    assign n4395 = n3050 ? encrypted_data_buf[1161] : n4387;   // modexp_top.v(481)
    assign n4396 = n3050 ? encrypted_data_buf[1160] : n4388;   // modexp_top.v(481)
    assign n4397 = n3044 ? encrypted_data_buf[1159] : n4389;   // modexp_top.v(481)
    assign n4398 = n3044 ? encrypted_data_buf[1158] : n4390;   // modexp_top.v(481)
    assign n4399 = n3044 ? encrypted_data_buf[1157] : n4391;   // modexp_top.v(481)
    assign n4400 = n3044 ? encrypted_data_buf[1156] : n4392;   // modexp_top.v(481)
    assign n4401 = n3044 ? encrypted_data_buf[1155] : n4393;   // modexp_top.v(481)
    assign n4402 = n3044 ? encrypted_data_buf[1154] : n4394;   // modexp_top.v(481)
    assign n4403 = n3044 ? encrypted_data_buf[1153] : n4395;   // modexp_top.v(481)
    assign n4404 = n3044 ? encrypted_data_buf[1152] : n4396;   // modexp_top.v(481)
    assign n4405 = n3037 ? encrypted_data_buf[1151] : n4397;   // modexp_top.v(481)
    assign n4406 = n3037 ? encrypted_data_buf[1150] : n4398;   // modexp_top.v(481)
    assign n4407 = n3037 ? encrypted_data_buf[1149] : n4399;   // modexp_top.v(481)
    assign n4408 = n3037 ? encrypted_data_buf[1148] : n4400;   // modexp_top.v(481)
    assign n4409 = n3037 ? encrypted_data_buf[1147] : n4401;   // modexp_top.v(481)
    assign n4410 = n3037 ? encrypted_data_buf[1146] : n4402;   // modexp_top.v(481)
    assign n4411 = n3037 ? encrypted_data_buf[1145] : n4403;   // modexp_top.v(481)
    assign n4412 = n3037 ? encrypted_data_buf[1144] : n4404;   // modexp_top.v(481)
    assign n4413 = n3033 ? encrypted_data_buf[1143] : n4405;   // modexp_top.v(481)
    assign n4414 = n3033 ? encrypted_data_buf[1142] : n4406;   // modexp_top.v(481)
    assign n4415 = n3033 ? encrypted_data_buf[1141] : n4407;   // modexp_top.v(481)
    assign n4416 = n3033 ? encrypted_data_buf[1140] : n4408;   // modexp_top.v(481)
    assign n4417 = n3033 ? encrypted_data_buf[1139] : n4409;   // modexp_top.v(481)
    assign n4418 = n3033 ? encrypted_data_buf[1138] : n4410;   // modexp_top.v(481)
    assign n4419 = n3033 ? encrypted_data_buf[1137] : n4411;   // modexp_top.v(481)
    assign n4420 = n3033 ? encrypted_data_buf[1136] : n4412;   // modexp_top.v(481)
    assign n4421 = n3028 ? encrypted_data_buf[1135] : n4413;   // modexp_top.v(481)
    assign n4422 = n3028 ? encrypted_data_buf[1134] : n4414;   // modexp_top.v(481)
    assign n4423 = n3028 ? encrypted_data_buf[1133] : n4415;   // modexp_top.v(481)
    assign n4424 = n3028 ? encrypted_data_buf[1132] : n4416;   // modexp_top.v(481)
    assign n4425 = n3028 ? encrypted_data_buf[1131] : n4417;   // modexp_top.v(481)
    assign n4426 = n3028 ? encrypted_data_buf[1130] : n4418;   // modexp_top.v(481)
    assign n4427 = n3028 ? encrypted_data_buf[1129] : n4419;   // modexp_top.v(481)
    assign n4428 = n3028 ? encrypted_data_buf[1128] : n4420;   // modexp_top.v(481)
    assign n4429 = n3023 ? encrypted_data_buf[1127] : n4421;   // modexp_top.v(481)
    assign n4430 = n3023 ? encrypted_data_buf[1126] : n4422;   // modexp_top.v(481)
    assign n4431 = n3023 ? encrypted_data_buf[1125] : n4423;   // modexp_top.v(481)
    assign n4432 = n3023 ? encrypted_data_buf[1124] : n4424;   // modexp_top.v(481)
    assign n4433 = n3023 ? encrypted_data_buf[1123] : n4425;   // modexp_top.v(481)
    assign n4434 = n3023 ? encrypted_data_buf[1122] : n4426;   // modexp_top.v(481)
    assign n4435 = n3023 ? encrypted_data_buf[1121] : n4427;   // modexp_top.v(481)
    assign n4436 = n3023 ? encrypted_data_buf[1120] : n4428;   // modexp_top.v(481)
    assign n4437 = n3017 ? encrypted_data_buf[1119] : n4429;   // modexp_top.v(481)
    assign n4438 = n3017 ? encrypted_data_buf[1118] : n4430;   // modexp_top.v(481)
    assign n4439 = n3017 ? encrypted_data_buf[1117] : n4431;   // modexp_top.v(481)
    assign n4440 = n3017 ? encrypted_data_buf[1116] : n4432;   // modexp_top.v(481)
    assign n4441 = n3017 ? encrypted_data_buf[1115] : n4433;   // modexp_top.v(481)
    assign n4442 = n3017 ? encrypted_data_buf[1114] : n4434;   // modexp_top.v(481)
    assign n4443 = n3017 ? encrypted_data_buf[1113] : n4435;   // modexp_top.v(481)
    assign n4444 = n3017 ? encrypted_data_buf[1112] : n4436;   // modexp_top.v(481)
    assign n4445 = n3012 ? encrypted_data_buf[1111] : n4437;   // modexp_top.v(481)
    assign n4446 = n3012 ? encrypted_data_buf[1110] : n4438;   // modexp_top.v(481)
    assign n4447 = n3012 ? encrypted_data_buf[1109] : n4439;   // modexp_top.v(481)
    assign n4448 = n3012 ? encrypted_data_buf[1108] : n4440;   // modexp_top.v(481)
    assign n4449 = n3012 ? encrypted_data_buf[1107] : n4441;   // modexp_top.v(481)
    assign n4450 = n3012 ? encrypted_data_buf[1106] : n4442;   // modexp_top.v(481)
    assign n4451 = n3012 ? encrypted_data_buf[1105] : n4443;   // modexp_top.v(481)
    assign n4452 = n3012 ? encrypted_data_buf[1104] : n4444;   // modexp_top.v(481)
    assign n4453 = n3006 ? encrypted_data_buf[1103] : n4445;   // modexp_top.v(481)
    assign n4454 = n3006 ? encrypted_data_buf[1102] : n4446;   // modexp_top.v(481)
    assign n4455 = n3006 ? encrypted_data_buf[1101] : n4447;   // modexp_top.v(481)
    assign n4456 = n3006 ? encrypted_data_buf[1100] : n4448;   // modexp_top.v(481)
    assign n4457 = n3006 ? encrypted_data_buf[1099] : n4449;   // modexp_top.v(481)
    assign n4458 = n3006 ? encrypted_data_buf[1098] : n4450;   // modexp_top.v(481)
    assign n4459 = n3006 ? encrypted_data_buf[1097] : n4451;   // modexp_top.v(481)
    assign n4460 = n3006 ? encrypted_data_buf[1096] : n4452;   // modexp_top.v(481)
    assign n4461 = n3000 ? encrypted_data_buf[1095] : n4453;   // modexp_top.v(481)
    assign n4462 = n3000 ? encrypted_data_buf[1094] : n4454;   // modexp_top.v(481)
    assign n4463 = n3000 ? encrypted_data_buf[1093] : n4455;   // modexp_top.v(481)
    assign n4464 = n3000 ? encrypted_data_buf[1092] : n4456;   // modexp_top.v(481)
    assign n4465 = n3000 ? encrypted_data_buf[1091] : n4457;   // modexp_top.v(481)
    assign n4466 = n3000 ? encrypted_data_buf[1090] : n4458;   // modexp_top.v(481)
    assign n4467 = n3000 ? encrypted_data_buf[1089] : n4459;   // modexp_top.v(481)
    assign n4468 = n3000 ? encrypted_data_buf[1088] : n4460;   // modexp_top.v(481)
    assign n4469 = n2993 ? encrypted_data_buf[1087] : n4461;   // modexp_top.v(481)
    assign n4470 = n2993 ? encrypted_data_buf[1086] : n4462;   // modexp_top.v(481)
    assign n4471 = n2993 ? encrypted_data_buf[1085] : n4463;   // modexp_top.v(481)
    assign n4472 = n2993 ? encrypted_data_buf[1084] : n4464;   // modexp_top.v(481)
    assign n4473 = n2993 ? encrypted_data_buf[1083] : n4465;   // modexp_top.v(481)
    assign n4474 = n2993 ? encrypted_data_buf[1082] : n4466;   // modexp_top.v(481)
    assign n4475 = n2993 ? encrypted_data_buf[1081] : n4467;   // modexp_top.v(481)
    assign n4476 = n2993 ? encrypted_data_buf[1080] : n4468;   // modexp_top.v(481)
    assign n4477 = n2988 ? encrypted_data_buf[1079] : n4469;   // modexp_top.v(481)
    assign n4478 = n2988 ? encrypted_data_buf[1078] : n4470;   // modexp_top.v(481)
    assign n4479 = n2988 ? encrypted_data_buf[1077] : n4471;   // modexp_top.v(481)
    assign n4480 = n2988 ? encrypted_data_buf[1076] : n4472;   // modexp_top.v(481)
    assign n4481 = n2988 ? encrypted_data_buf[1075] : n4473;   // modexp_top.v(481)
    assign n4482 = n2988 ? encrypted_data_buf[1074] : n4474;   // modexp_top.v(481)
    assign n4483 = n2988 ? encrypted_data_buf[1073] : n4475;   // modexp_top.v(481)
    assign n4484 = n2988 ? encrypted_data_buf[1072] : n4476;   // modexp_top.v(481)
    assign n4485 = n2982 ? encrypted_data_buf[1071] : n4477;   // modexp_top.v(481)
    assign n4486 = n2982 ? encrypted_data_buf[1070] : n4478;   // modexp_top.v(481)
    assign n4487 = n2982 ? encrypted_data_buf[1069] : n4479;   // modexp_top.v(481)
    assign n4488 = n2982 ? encrypted_data_buf[1068] : n4480;   // modexp_top.v(481)
    assign n4489 = n2982 ? encrypted_data_buf[1067] : n4481;   // modexp_top.v(481)
    assign n4490 = n2982 ? encrypted_data_buf[1066] : n4482;   // modexp_top.v(481)
    assign n4491 = n2982 ? encrypted_data_buf[1065] : n4483;   // modexp_top.v(481)
    assign n4492 = n2982 ? encrypted_data_buf[1064] : n4484;   // modexp_top.v(481)
    assign n4493 = n2976 ? encrypted_data_buf[1063] : n4485;   // modexp_top.v(481)
    assign n4494 = n2976 ? encrypted_data_buf[1062] : n4486;   // modexp_top.v(481)
    assign n4495 = n2976 ? encrypted_data_buf[1061] : n4487;   // modexp_top.v(481)
    assign n4496 = n2976 ? encrypted_data_buf[1060] : n4488;   // modexp_top.v(481)
    assign n4497 = n2976 ? encrypted_data_buf[1059] : n4489;   // modexp_top.v(481)
    assign n4498 = n2976 ? encrypted_data_buf[1058] : n4490;   // modexp_top.v(481)
    assign n4499 = n2976 ? encrypted_data_buf[1057] : n4491;   // modexp_top.v(481)
    assign n4500 = n2976 ? encrypted_data_buf[1056] : n4492;   // modexp_top.v(481)
    assign n4501 = n2969 ? encrypted_data_buf[1055] : n4493;   // modexp_top.v(481)
    assign n4502 = n2969 ? encrypted_data_buf[1054] : n4494;   // modexp_top.v(481)
    assign n4503 = n2969 ? encrypted_data_buf[1053] : n4495;   // modexp_top.v(481)
    assign n4504 = n2969 ? encrypted_data_buf[1052] : n4496;   // modexp_top.v(481)
    assign n4505 = n2969 ? encrypted_data_buf[1051] : n4497;   // modexp_top.v(481)
    assign n4506 = n2969 ? encrypted_data_buf[1050] : n4498;   // modexp_top.v(481)
    assign n4507 = n2969 ? encrypted_data_buf[1049] : n4499;   // modexp_top.v(481)
    assign n4508 = n2969 ? encrypted_data_buf[1048] : n4500;   // modexp_top.v(481)
    assign n4509 = n2963 ? encrypted_data_buf[1047] : n4501;   // modexp_top.v(481)
    assign n4510 = n2963 ? encrypted_data_buf[1046] : n4502;   // modexp_top.v(481)
    assign n4511 = n2963 ? encrypted_data_buf[1045] : n4503;   // modexp_top.v(481)
    assign n4512 = n2963 ? encrypted_data_buf[1044] : n4504;   // modexp_top.v(481)
    assign n4513 = n2963 ? encrypted_data_buf[1043] : n4505;   // modexp_top.v(481)
    assign n4514 = n2963 ? encrypted_data_buf[1042] : n4506;   // modexp_top.v(481)
    assign n4515 = n2963 ? encrypted_data_buf[1041] : n4507;   // modexp_top.v(481)
    assign n4516 = n2963 ? encrypted_data_buf[1040] : n4508;   // modexp_top.v(481)
    assign n4517 = n2956 ? encrypted_data_buf[1039] : n4509;   // modexp_top.v(481)
    assign n4518 = n2956 ? encrypted_data_buf[1038] : n4510;   // modexp_top.v(481)
    assign n4519 = n2956 ? encrypted_data_buf[1037] : n4511;   // modexp_top.v(481)
    assign n4520 = n2956 ? encrypted_data_buf[1036] : n4512;   // modexp_top.v(481)
    assign n4521 = n2956 ? encrypted_data_buf[1035] : n4513;   // modexp_top.v(481)
    assign n4522 = n2956 ? encrypted_data_buf[1034] : n4514;   // modexp_top.v(481)
    assign n4523 = n2956 ? encrypted_data_buf[1033] : n4515;   // modexp_top.v(481)
    assign n4524 = n2956 ? encrypted_data_buf[1032] : n4516;   // modexp_top.v(481)
    assign n4525 = n2949 ? encrypted_data_buf[1031] : n4517;   // modexp_top.v(481)
    assign n4526 = n2949 ? encrypted_data_buf[1030] : n4518;   // modexp_top.v(481)
    assign n4527 = n2949 ? encrypted_data_buf[1029] : n4519;   // modexp_top.v(481)
    assign n4528 = n2949 ? encrypted_data_buf[1028] : n4520;   // modexp_top.v(481)
    assign n4529 = n2949 ? encrypted_data_buf[1027] : n4521;   // modexp_top.v(481)
    assign n4530 = n2949 ? encrypted_data_buf[1026] : n4522;   // modexp_top.v(481)
    assign n4531 = n2949 ? encrypted_data_buf[1025] : n4523;   // modexp_top.v(481)
    assign n4532 = n2949 ? encrypted_data_buf[1024] : n4524;   // modexp_top.v(481)
    assign n4533 = n2941 ? encrypted_data_buf[1023] : n4525;   // modexp_top.v(481)
    assign n4534 = n2941 ? encrypted_data_buf[1022] : n4526;   // modexp_top.v(481)
    assign n4535 = n2941 ? encrypted_data_buf[1021] : n4527;   // modexp_top.v(481)
    assign n4536 = n2941 ? encrypted_data_buf[1020] : n4528;   // modexp_top.v(481)
    assign n4537 = n2941 ? encrypted_data_buf[1019] : n4529;   // modexp_top.v(481)
    assign n4538 = n2941 ? encrypted_data_buf[1018] : n4530;   // modexp_top.v(481)
    assign n4539 = n2941 ? encrypted_data_buf[1017] : n4531;   // modexp_top.v(481)
    assign n4540 = n2941 ? encrypted_data_buf[1016] : n4532;   // modexp_top.v(481)
    assign n4541 = n2939 ? encrypted_data_buf[1015] : n4533;   // modexp_top.v(481)
    assign n4542 = n2939 ? encrypted_data_buf[1014] : n4534;   // modexp_top.v(481)
    assign n4543 = n2939 ? encrypted_data_buf[1013] : n4535;   // modexp_top.v(481)
    assign n4544 = n2939 ? encrypted_data_buf[1012] : n4536;   // modexp_top.v(481)
    assign n4545 = n2939 ? encrypted_data_buf[1011] : n4537;   // modexp_top.v(481)
    assign n4546 = n2939 ? encrypted_data_buf[1010] : n4538;   // modexp_top.v(481)
    assign n4547 = n2939 ? encrypted_data_buf[1009] : n4539;   // modexp_top.v(481)
    assign n4548 = n2939 ? encrypted_data_buf[1008] : n4540;   // modexp_top.v(481)
    assign n4549 = n2936 ? encrypted_data_buf[1007] : n4541;   // modexp_top.v(481)
    assign n4550 = n2936 ? encrypted_data_buf[1006] : n4542;   // modexp_top.v(481)
    assign n4551 = n2936 ? encrypted_data_buf[1005] : n4543;   // modexp_top.v(481)
    assign n4552 = n2936 ? encrypted_data_buf[1004] : n4544;   // modexp_top.v(481)
    assign n4553 = n2936 ? encrypted_data_buf[1003] : n4545;   // modexp_top.v(481)
    assign n4554 = n2936 ? encrypted_data_buf[1002] : n4546;   // modexp_top.v(481)
    assign n4555 = n2936 ? encrypted_data_buf[1001] : n4547;   // modexp_top.v(481)
    assign n4556 = n2936 ? encrypted_data_buf[1000] : n4548;   // modexp_top.v(481)
    assign n4557 = n2933 ? encrypted_data_buf[999] : n4549;   // modexp_top.v(481)
    assign n4558 = n2933 ? encrypted_data_buf[998] : n4550;   // modexp_top.v(481)
    assign n4559 = n2933 ? encrypted_data_buf[997] : n4551;   // modexp_top.v(481)
    assign n4560 = n2933 ? encrypted_data_buf[996] : n4552;   // modexp_top.v(481)
    assign n4561 = n2933 ? encrypted_data_buf[995] : n4553;   // modexp_top.v(481)
    assign n4562 = n2933 ? encrypted_data_buf[994] : n4554;   // modexp_top.v(481)
    assign n4563 = n2933 ? encrypted_data_buf[993] : n4555;   // modexp_top.v(481)
    assign n4564 = n2933 ? encrypted_data_buf[992] : n4556;   // modexp_top.v(481)
    assign n4565 = n2929 ? encrypted_data_buf[991] : n4557;   // modexp_top.v(481)
    assign n4566 = n2929 ? encrypted_data_buf[990] : n4558;   // modexp_top.v(481)
    assign n4567 = n2929 ? encrypted_data_buf[989] : n4559;   // modexp_top.v(481)
    assign n4568 = n2929 ? encrypted_data_buf[988] : n4560;   // modexp_top.v(481)
    assign n4569 = n2929 ? encrypted_data_buf[987] : n4561;   // modexp_top.v(481)
    assign n4570 = n2929 ? encrypted_data_buf[986] : n4562;   // modexp_top.v(481)
    assign n4571 = n2929 ? encrypted_data_buf[985] : n4563;   // modexp_top.v(481)
    assign n4572 = n2929 ? encrypted_data_buf[984] : n4564;   // modexp_top.v(481)
    assign n4573 = n2926 ? encrypted_data_buf[983] : n4565;   // modexp_top.v(481)
    assign n4574 = n2926 ? encrypted_data_buf[982] : n4566;   // modexp_top.v(481)
    assign n4575 = n2926 ? encrypted_data_buf[981] : n4567;   // modexp_top.v(481)
    assign n4576 = n2926 ? encrypted_data_buf[980] : n4568;   // modexp_top.v(481)
    assign n4577 = n2926 ? encrypted_data_buf[979] : n4569;   // modexp_top.v(481)
    assign n4578 = n2926 ? encrypted_data_buf[978] : n4570;   // modexp_top.v(481)
    assign n4579 = n2926 ? encrypted_data_buf[977] : n4571;   // modexp_top.v(481)
    assign n4580 = n2926 ? encrypted_data_buf[976] : n4572;   // modexp_top.v(481)
    assign n4581 = n2922 ? encrypted_data_buf[975] : n4573;   // modexp_top.v(481)
    assign n4582 = n2922 ? encrypted_data_buf[974] : n4574;   // modexp_top.v(481)
    assign n4583 = n2922 ? encrypted_data_buf[973] : n4575;   // modexp_top.v(481)
    assign n4584 = n2922 ? encrypted_data_buf[972] : n4576;   // modexp_top.v(481)
    assign n4585 = n2922 ? encrypted_data_buf[971] : n4577;   // modexp_top.v(481)
    assign n4586 = n2922 ? encrypted_data_buf[970] : n4578;   // modexp_top.v(481)
    assign n4587 = n2922 ? encrypted_data_buf[969] : n4579;   // modexp_top.v(481)
    assign n4588 = n2922 ? encrypted_data_buf[968] : n4580;   // modexp_top.v(481)
    assign n4589 = n2918 ? encrypted_data_buf[967] : n4581;   // modexp_top.v(481)
    assign n4590 = n2918 ? encrypted_data_buf[966] : n4582;   // modexp_top.v(481)
    assign n4591 = n2918 ? encrypted_data_buf[965] : n4583;   // modexp_top.v(481)
    assign n4592 = n2918 ? encrypted_data_buf[964] : n4584;   // modexp_top.v(481)
    assign n4593 = n2918 ? encrypted_data_buf[963] : n4585;   // modexp_top.v(481)
    assign n4594 = n2918 ? encrypted_data_buf[962] : n4586;   // modexp_top.v(481)
    assign n4595 = n2918 ? encrypted_data_buf[961] : n4587;   // modexp_top.v(481)
    assign n4596 = n2918 ? encrypted_data_buf[960] : n4588;   // modexp_top.v(481)
    assign n4597 = n2913 ? encrypted_data_buf[959] : n4589;   // modexp_top.v(481)
    assign n4598 = n2913 ? encrypted_data_buf[958] : n4590;   // modexp_top.v(481)
    assign n4599 = n2913 ? encrypted_data_buf[957] : n4591;   // modexp_top.v(481)
    assign n4600 = n2913 ? encrypted_data_buf[956] : n4592;   // modexp_top.v(481)
    assign n4601 = n2913 ? encrypted_data_buf[955] : n4593;   // modexp_top.v(481)
    assign n4602 = n2913 ? encrypted_data_buf[954] : n4594;   // modexp_top.v(481)
    assign n4603 = n2913 ? encrypted_data_buf[953] : n4595;   // modexp_top.v(481)
    assign n4604 = n2913 ? encrypted_data_buf[952] : n4596;   // modexp_top.v(481)
    assign n4605 = n2910 ? encrypted_data_buf[951] : n4597;   // modexp_top.v(481)
    assign n4606 = n2910 ? encrypted_data_buf[950] : n4598;   // modexp_top.v(481)
    assign n4607 = n2910 ? encrypted_data_buf[949] : n4599;   // modexp_top.v(481)
    assign n4608 = n2910 ? encrypted_data_buf[948] : n4600;   // modexp_top.v(481)
    assign n4609 = n2910 ? encrypted_data_buf[947] : n4601;   // modexp_top.v(481)
    assign n4610 = n2910 ? encrypted_data_buf[946] : n4602;   // modexp_top.v(481)
    assign n4611 = n2910 ? encrypted_data_buf[945] : n4603;   // modexp_top.v(481)
    assign n4612 = n2910 ? encrypted_data_buf[944] : n4604;   // modexp_top.v(481)
    assign n4613 = n2906 ? encrypted_data_buf[943] : n4605;   // modexp_top.v(481)
    assign n4614 = n2906 ? encrypted_data_buf[942] : n4606;   // modexp_top.v(481)
    assign n4615 = n2906 ? encrypted_data_buf[941] : n4607;   // modexp_top.v(481)
    assign n4616 = n2906 ? encrypted_data_buf[940] : n4608;   // modexp_top.v(481)
    assign n4617 = n2906 ? encrypted_data_buf[939] : n4609;   // modexp_top.v(481)
    assign n4618 = n2906 ? encrypted_data_buf[938] : n4610;   // modexp_top.v(481)
    assign n4619 = n2906 ? encrypted_data_buf[937] : n4611;   // modexp_top.v(481)
    assign n4620 = n2906 ? encrypted_data_buf[936] : n4612;   // modexp_top.v(481)
    assign n4621 = n2902 ? encrypted_data_buf[935] : n4613;   // modexp_top.v(481)
    assign n4622 = n2902 ? encrypted_data_buf[934] : n4614;   // modexp_top.v(481)
    assign n4623 = n2902 ? encrypted_data_buf[933] : n4615;   // modexp_top.v(481)
    assign n4624 = n2902 ? encrypted_data_buf[932] : n4616;   // modexp_top.v(481)
    assign n4625 = n2902 ? encrypted_data_buf[931] : n4617;   // modexp_top.v(481)
    assign n4626 = n2902 ? encrypted_data_buf[930] : n4618;   // modexp_top.v(481)
    assign n4627 = n2902 ? encrypted_data_buf[929] : n4619;   // modexp_top.v(481)
    assign n4628 = n2902 ? encrypted_data_buf[928] : n4620;   // modexp_top.v(481)
    assign n4629 = n2897 ? encrypted_data_buf[927] : n4621;   // modexp_top.v(481)
    assign n4630 = n2897 ? encrypted_data_buf[926] : n4622;   // modexp_top.v(481)
    assign n4631 = n2897 ? encrypted_data_buf[925] : n4623;   // modexp_top.v(481)
    assign n4632 = n2897 ? encrypted_data_buf[924] : n4624;   // modexp_top.v(481)
    assign n4633 = n2897 ? encrypted_data_buf[923] : n4625;   // modexp_top.v(481)
    assign n4634 = n2897 ? encrypted_data_buf[922] : n4626;   // modexp_top.v(481)
    assign n4635 = n2897 ? encrypted_data_buf[921] : n4627;   // modexp_top.v(481)
    assign n4636 = n2897 ? encrypted_data_buf[920] : n4628;   // modexp_top.v(481)
    assign n4637 = n2893 ? encrypted_data_buf[919] : n4629;   // modexp_top.v(481)
    assign n4638 = n2893 ? encrypted_data_buf[918] : n4630;   // modexp_top.v(481)
    assign n4639 = n2893 ? encrypted_data_buf[917] : n4631;   // modexp_top.v(481)
    assign n4640 = n2893 ? encrypted_data_buf[916] : n4632;   // modexp_top.v(481)
    assign n4641 = n2893 ? encrypted_data_buf[915] : n4633;   // modexp_top.v(481)
    assign n4642 = n2893 ? encrypted_data_buf[914] : n4634;   // modexp_top.v(481)
    assign n4643 = n2893 ? encrypted_data_buf[913] : n4635;   // modexp_top.v(481)
    assign n4644 = n2893 ? encrypted_data_buf[912] : n4636;   // modexp_top.v(481)
    assign n4645 = n2888 ? encrypted_data_buf[911] : n4637;   // modexp_top.v(481)
    assign n4646 = n2888 ? encrypted_data_buf[910] : n4638;   // modexp_top.v(481)
    assign n4647 = n2888 ? encrypted_data_buf[909] : n4639;   // modexp_top.v(481)
    assign n4648 = n2888 ? encrypted_data_buf[908] : n4640;   // modexp_top.v(481)
    assign n4649 = n2888 ? encrypted_data_buf[907] : n4641;   // modexp_top.v(481)
    assign n4650 = n2888 ? encrypted_data_buf[906] : n4642;   // modexp_top.v(481)
    assign n4651 = n2888 ? encrypted_data_buf[905] : n4643;   // modexp_top.v(481)
    assign n4652 = n2888 ? encrypted_data_buf[904] : n4644;   // modexp_top.v(481)
    assign n4653 = n2883 ? encrypted_data_buf[903] : n4645;   // modexp_top.v(481)
    assign n4654 = n2883 ? encrypted_data_buf[902] : n4646;   // modexp_top.v(481)
    assign n4655 = n2883 ? encrypted_data_buf[901] : n4647;   // modexp_top.v(481)
    assign n4656 = n2883 ? encrypted_data_buf[900] : n4648;   // modexp_top.v(481)
    assign n4657 = n2883 ? encrypted_data_buf[899] : n4649;   // modexp_top.v(481)
    assign n4658 = n2883 ? encrypted_data_buf[898] : n4650;   // modexp_top.v(481)
    assign n4659 = n2883 ? encrypted_data_buf[897] : n4651;   // modexp_top.v(481)
    assign n4660 = n2883 ? encrypted_data_buf[896] : n4652;   // modexp_top.v(481)
    assign n4661 = n2877 ? encrypted_data_buf[895] : n4653;   // modexp_top.v(481)
    assign n4662 = n2877 ? encrypted_data_buf[894] : n4654;   // modexp_top.v(481)
    assign n4663 = n2877 ? encrypted_data_buf[893] : n4655;   // modexp_top.v(481)
    assign n4664 = n2877 ? encrypted_data_buf[892] : n4656;   // modexp_top.v(481)
    assign n4665 = n2877 ? encrypted_data_buf[891] : n4657;   // modexp_top.v(481)
    assign n4666 = n2877 ? encrypted_data_buf[890] : n4658;   // modexp_top.v(481)
    assign n4667 = n2877 ? encrypted_data_buf[889] : n4659;   // modexp_top.v(481)
    assign n4668 = n2877 ? encrypted_data_buf[888] : n4660;   // modexp_top.v(481)
    assign n4669 = n2874 ? encrypted_data_buf[887] : n4661;   // modexp_top.v(481)
    assign n4670 = n2874 ? encrypted_data_buf[886] : n4662;   // modexp_top.v(481)
    assign n4671 = n2874 ? encrypted_data_buf[885] : n4663;   // modexp_top.v(481)
    assign n4672 = n2874 ? encrypted_data_buf[884] : n4664;   // modexp_top.v(481)
    assign n4673 = n2874 ? encrypted_data_buf[883] : n4665;   // modexp_top.v(481)
    assign n4674 = n2874 ? encrypted_data_buf[882] : n4666;   // modexp_top.v(481)
    assign n4675 = n2874 ? encrypted_data_buf[881] : n4667;   // modexp_top.v(481)
    assign n4676 = n2874 ? encrypted_data_buf[880] : n4668;   // modexp_top.v(481)
    assign n4677 = n2870 ? encrypted_data_buf[879] : n4669;   // modexp_top.v(481)
    assign n4678 = n2870 ? encrypted_data_buf[878] : n4670;   // modexp_top.v(481)
    assign n4679 = n2870 ? encrypted_data_buf[877] : n4671;   // modexp_top.v(481)
    assign n4680 = n2870 ? encrypted_data_buf[876] : n4672;   // modexp_top.v(481)
    assign n4681 = n2870 ? encrypted_data_buf[875] : n4673;   // modexp_top.v(481)
    assign n4682 = n2870 ? encrypted_data_buf[874] : n4674;   // modexp_top.v(481)
    assign n4683 = n2870 ? encrypted_data_buf[873] : n4675;   // modexp_top.v(481)
    assign n4684 = n2870 ? encrypted_data_buf[872] : n4676;   // modexp_top.v(481)
    assign n4685 = n2866 ? encrypted_data_buf[871] : n4677;   // modexp_top.v(481)
    assign n4686 = n2866 ? encrypted_data_buf[870] : n4678;   // modexp_top.v(481)
    assign n4687 = n2866 ? encrypted_data_buf[869] : n4679;   // modexp_top.v(481)
    assign n4688 = n2866 ? encrypted_data_buf[868] : n4680;   // modexp_top.v(481)
    assign n4689 = n2866 ? encrypted_data_buf[867] : n4681;   // modexp_top.v(481)
    assign n4690 = n2866 ? encrypted_data_buf[866] : n4682;   // modexp_top.v(481)
    assign n4691 = n2866 ? encrypted_data_buf[865] : n4683;   // modexp_top.v(481)
    assign n4692 = n2866 ? encrypted_data_buf[864] : n4684;   // modexp_top.v(481)
    assign n4693 = n2861 ? encrypted_data_buf[863] : n4685;   // modexp_top.v(481)
    assign n4694 = n2861 ? encrypted_data_buf[862] : n4686;   // modexp_top.v(481)
    assign n4695 = n2861 ? encrypted_data_buf[861] : n4687;   // modexp_top.v(481)
    assign n4696 = n2861 ? encrypted_data_buf[860] : n4688;   // modexp_top.v(481)
    assign n4697 = n2861 ? encrypted_data_buf[859] : n4689;   // modexp_top.v(481)
    assign n4698 = n2861 ? encrypted_data_buf[858] : n4690;   // modexp_top.v(481)
    assign n4699 = n2861 ? encrypted_data_buf[857] : n4691;   // modexp_top.v(481)
    assign n4700 = n2861 ? encrypted_data_buf[856] : n4692;   // modexp_top.v(481)
    assign n4701 = n2857 ? encrypted_data_buf[855] : n4693;   // modexp_top.v(481)
    assign n4702 = n2857 ? encrypted_data_buf[854] : n4694;   // modexp_top.v(481)
    assign n4703 = n2857 ? encrypted_data_buf[853] : n4695;   // modexp_top.v(481)
    assign n4704 = n2857 ? encrypted_data_buf[852] : n4696;   // modexp_top.v(481)
    assign n4705 = n2857 ? encrypted_data_buf[851] : n4697;   // modexp_top.v(481)
    assign n4706 = n2857 ? encrypted_data_buf[850] : n4698;   // modexp_top.v(481)
    assign n4707 = n2857 ? encrypted_data_buf[849] : n4699;   // modexp_top.v(481)
    assign n4708 = n2857 ? encrypted_data_buf[848] : n4700;   // modexp_top.v(481)
    assign n4709 = n2852 ? encrypted_data_buf[847] : n4701;   // modexp_top.v(481)
    assign n4710 = n2852 ? encrypted_data_buf[846] : n4702;   // modexp_top.v(481)
    assign n4711 = n2852 ? encrypted_data_buf[845] : n4703;   // modexp_top.v(481)
    assign n4712 = n2852 ? encrypted_data_buf[844] : n4704;   // modexp_top.v(481)
    assign n4713 = n2852 ? encrypted_data_buf[843] : n4705;   // modexp_top.v(481)
    assign n4714 = n2852 ? encrypted_data_buf[842] : n4706;   // modexp_top.v(481)
    assign n4715 = n2852 ? encrypted_data_buf[841] : n4707;   // modexp_top.v(481)
    assign n4716 = n2852 ? encrypted_data_buf[840] : n4708;   // modexp_top.v(481)
    assign n4717 = n2847 ? encrypted_data_buf[839] : n4709;   // modexp_top.v(481)
    assign n4718 = n2847 ? encrypted_data_buf[838] : n4710;   // modexp_top.v(481)
    assign n4719 = n2847 ? encrypted_data_buf[837] : n4711;   // modexp_top.v(481)
    assign n4720 = n2847 ? encrypted_data_buf[836] : n4712;   // modexp_top.v(481)
    assign n4721 = n2847 ? encrypted_data_buf[835] : n4713;   // modexp_top.v(481)
    assign n4722 = n2847 ? encrypted_data_buf[834] : n4714;   // modexp_top.v(481)
    assign n4723 = n2847 ? encrypted_data_buf[833] : n4715;   // modexp_top.v(481)
    assign n4724 = n2847 ? encrypted_data_buf[832] : n4716;   // modexp_top.v(481)
    assign n4725 = n2841 ? encrypted_data_buf[831] : n4717;   // modexp_top.v(481)
    assign n4726 = n2841 ? encrypted_data_buf[830] : n4718;   // modexp_top.v(481)
    assign n4727 = n2841 ? encrypted_data_buf[829] : n4719;   // modexp_top.v(481)
    assign n4728 = n2841 ? encrypted_data_buf[828] : n4720;   // modexp_top.v(481)
    assign n4729 = n2841 ? encrypted_data_buf[827] : n4721;   // modexp_top.v(481)
    assign n4730 = n2841 ? encrypted_data_buf[826] : n4722;   // modexp_top.v(481)
    assign n4731 = n2841 ? encrypted_data_buf[825] : n4723;   // modexp_top.v(481)
    assign n4732 = n2841 ? encrypted_data_buf[824] : n4724;   // modexp_top.v(481)
    assign n4733 = n2837 ? encrypted_data_buf[823] : n4725;   // modexp_top.v(481)
    assign n4734 = n2837 ? encrypted_data_buf[822] : n4726;   // modexp_top.v(481)
    assign n4735 = n2837 ? encrypted_data_buf[821] : n4727;   // modexp_top.v(481)
    assign n4736 = n2837 ? encrypted_data_buf[820] : n4728;   // modexp_top.v(481)
    assign n4737 = n2837 ? encrypted_data_buf[819] : n4729;   // modexp_top.v(481)
    assign n4738 = n2837 ? encrypted_data_buf[818] : n4730;   // modexp_top.v(481)
    assign n4739 = n2837 ? encrypted_data_buf[817] : n4731;   // modexp_top.v(481)
    assign n4740 = n2837 ? encrypted_data_buf[816] : n4732;   // modexp_top.v(481)
    assign n4741 = n2832 ? encrypted_data_buf[815] : n4733;   // modexp_top.v(481)
    assign n4742 = n2832 ? encrypted_data_buf[814] : n4734;   // modexp_top.v(481)
    assign n4743 = n2832 ? encrypted_data_buf[813] : n4735;   // modexp_top.v(481)
    assign n4744 = n2832 ? encrypted_data_buf[812] : n4736;   // modexp_top.v(481)
    assign n4745 = n2832 ? encrypted_data_buf[811] : n4737;   // modexp_top.v(481)
    assign n4746 = n2832 ? encrypted_data_buf[810] : n4738;   // modexp_top.v(481)
    assign n4747 = n2832 ? encrypted_data_buf[809] : n4739;   // modexp_top.v(481)
    assign n4748 = n2832 ? encrypted_data_buf[808] : n4740;   // modexp_top.v(481)
    assign n4749 = n2827 ? encrypted_data_buf[807] : n4741;   // modexp_top.v(481)
    assign n4750 = n2827 ? encrypted_data_buf[806] : n4742;   // modexp_top.v(481)
    assign n4751 = n2827 ? encrypted_data_buf[805] : n4743;   // modexp_top.v(481)
    assign n4752 = n2827 ? encrypted_data_buf[804] : n4744;   // modexp_top.v(481)
    assign n4753 = n2827 ? encrypted_data_buf[803] : n4745;   // modexp_top.v(481)
    assign n4754 = n2827 ? encrypted_data_buf[802] : n4746;   // modexp_top.v(481)
    assign n4755 = n2827 ? encrypted_data_buf[801] : n4747;   // modexp_top.v(481)
    assign n4756 = n2827 ? encrypted_data_buf[800] : n4748;   // modexp_top.v(481)
    assign n4757 = n2821 ? encrypted_data_buf[799] : n4749;   // modexp_top.v(481)
    assign n4758 = n2821 ? encrypted_data_buf[798] : n4750;   // modexp_top.v(481)
    assign n4759 = n2821 ? encrypted_data_buf[797] : n4751;   // modexp_top.v(481)
    assign n4760 = n2821 ? encrypted_data_buf[796] : n4752;   // modexp_top.v(481)
    assign n4761 = n2821 ? encrypted_data_buf[795] : n4753;   // modexp_top.v(481)
    assign n4762 = n2821 ? encrypted_data_buf[794] : n4754;   // modexp_top.v(481)
    assign n4763 = n2821 ? encrypted_data_buf[793] : n4755;   // modexp_top.v(481)
    assign n4764 = n2821 ? encrypted_data_buf[792] : n4756;   // modexp_top.v(481)
    assign n4765 = n2816 ? encrypted_data_buf[791] : n4757;   // modexp_top.v(481)
    assign n4766 = n2816 ? encrypted_data_buf[790] : n4758;   // modexp_top.v(481)
    assign n4767 = n2816 ? encrypted_data_buf[789] : n4759;   // modexp_top.v(481)
    assign n4768 = n2816 ? encrypted_data_buf[788] : n4760;   // modexp_top.v(481)
    assign n4769 = n2816 ? encrypted_data_buf[787] : n4761;   // modexp_top.v(481)
    assign n4770 = n2816 ? encrypted_data_buf[786] : n4762;   // modexp_top.v(481)
    assign n4771 = n2816 ? encrypted_data_buf[785] : n4763;   // modexp_top.v(481)
    assign n4772 = n2816 ? encrypted_data_buf[784] : n4764;   // modexp_top.v(481)
    assign n4773 = n2810 ? encrypted_data_buf[783] : n4765;   // modexp_top.v(481)
    assign n4774 = n2810 ? encrypted_data_buf[782] : n4766;   // modexp_top.v(481)
    assign n4775 = n2810 ? encrypted_data_buf[781] : n4767;   // modexp_top.v(481)
    assign n4776 = n2810 ? encrypted_data_buf[780] : n4768;   // modexp_top.v(481)
    assign n4777 = n2810 ? encrypted_data_buf[779] : n4769;   // modexp_top.v(481)
    assign n4778 = n2810 ? encrypted_data_buf[778] : n4770;   // modexp_top.v(481)
    assign n4779 = n2810 ? encrypted_data_buf[777] : n4771;   // modexp_top.v(481)
    assign n4780 = n2810 ? encrypted_data_buf[776] : n4772;   // modexp_top.v(481)
    assign n4781 = n2804 ? encrypted_data_buf[775] : n4773;   // modexp_top.v(481)
    assign n4782 = n2804 ? encrypted_data_buf[774] : n4774;   // modexp_top.v(481)
    assign n4783 = n2804 ? encrypted_data_buf[773] : n4775;   // modexp_top.v(481)
    assign n4784 = n2804 ? encrypted_data_buf[772] : n4776;   // modexp_top.v(481)
    assign n4785 = n2804 ? encrypted_data_buf[771] : n4777;   // modexp_top.v(481)
    assign n4786 = n2804 ? encrypted_data_buf[770] : n4778;   // modexp_top.v(481)
    assign n4787 = n2804 ? encrypted_data_buf[769] : n4779;   // modexp_top.v(481)
    assign n4788 = n2804 ? encrypted_data_buf[768] : n4780;   // modexp_top.v(481)
    assign n4789 = n2797 ? encrypted_data_buf[767] : n4781;   // modexp_top.v(481)
    assign n4790 = n2797 ? encrypted_data_buf[766] : n4782;   // modexp_top.v(481)
    assign n4791 = n2797 ? encrypted_data_buf[765] : n4783;   // modexp_top.v(481)
    assign n4792 = n2797 ? encrypted_data_buf[764] : n4784;   // modexp_top.v(481)
    assign n4793 = n2797 ? encrypted_data_buf[763] : n4785;   // modexp_top.v(481)
    assign n4794 = n2797 ? encrypted_data_buf[762] : n4786;   // modexp_top.v(481)
    assign n4795 = n2797 ? encrypted_data_buf[761] : n4787;   // modexp_top.v(481)
    assign n4796 = n2797 ? encrypted_data_buf[760] : n4788;   // modexp_top.v(481)
    assign n4797 = n2794 ? encrypted_data_buf[759] : n4789;   // modexp_top.v(481)
    assign n4798 = n2794 ? encrypted_data_buf[758] : n4790;   // modexp_top.v(481)
    assign n4799 = n2794 ? encrypted_data_buf[757] : n4791;   // modexp_top.v(481)
    assign n4800 = n2794 ? encrypted_data_buf[756] : n4792;   // modexp_top.v(481)
    assign n4801 = n2794 ? encrypted_data_buf[755] : n4793;   // modexp_top.v(481)
    assign n4802 = n2794 ? encrypted_data_buf[754] : n4794;   // modexp_top.v(481)
    assign n4803 = n2794 ? encrypted_data_buf[753] : n4795;   // modexp_top.v(481)
    assign n4804 = n2794 ? encrypted_data_buf[752] : n4796;   // modexp_top.v(481)
    assign n4805 = n2790 ? encrypted_data_buf[751] : n4797;   // modexp_top.v(481)
    assign n4806 = n2790 ? encrypted_data_buf[750] : n4798;   // modexp_top.v(481)
    assign n4807 = n2790 ? encrypted_data_buf[749] : n4799;   // modexp_top.v(481)
    assign n4808 = n2790 ? encrypted_data_buf[748] : n4800;   // modexp_top.v(481)
    assign n4809 = n2790 ? encrypted_data_buf[747] : n4801;   // modexp_top.v(481)
    assign n4810 = n2790 ? encrypted_data_buf[746] : n4802;   // modexp_top.v(481)
    assign n4811 = n2790 ? encrypted_data_buf[745] : n4803;   // modexp_top.v(481)
    assign n4812 = n2790 ? encrypted_data_buf[744] : n4804;   // modexp_top.v(481)
    assign n4813 = n2786 ? encrypted_data_buf[743] : n4805;   // modexp_top.v(481)
    assign n4814 = n2786 ? encrypted_data_buf[742] : n4806;   // modexp_top.v(481)
    assign n4815 = n2786 ? encrypted_data_buf[741] : n4807;   // modexp_top.v(481)
    assign n4816 = n2786 ? encrypted_data_buf[740] : n4808;   // modexp_top.v(481)
    assign n4817 = n2786 ? encrypted_data_buf[739] : n4809;   // modexp_top.v(481)
    assign n4818 = n2786 ? encrypted_data_buf[738] : n4810;   // modexp_top.v(481)
    assign n4819 = n2786 ? encrypted_data_buf[737] : n4811;   // modexp_top.v(481)
    assign n4820 = n2786 ? encrypted_data_buf[736] : n4812;   // modexp_top.v(481)
    assign n4821 = n2781 ? encrypted_data_buf[735] : n4813;   // modexp_top.v(481)
    assign n4822 = n2781 ? encrypted_data_buf[734] : n4814;   // modexp_top.v(481)
    assign n4823 = n2781 ? encrypted_data_buf[733] : n4815;   // modexp_top.v(481)
    assign n4824 = n2781 ? encrypted_data_buf[732] : n4816;   // modexp_top.v(481)
    assign n4825 = n2781 ? encrypted_data_buf[731] : n4817;   // modexp_top.v(481)
    assign n4826 = n2781 ? encrypted_data_buf[730] : n4818;   // modexp_top.v(481)
    assign n4827 = n2781 ? encrypted_data_buf[729] : n4819;   // modexp_top.v(481)
    assign n4828 = n2781 ? encrypted_data_buf[728] : n4820;   // modexp_top.v(481)
    assign n4829 = n2777 ? encrypted_data_buf[727] : n4821;   // modexp_top.v(481)
    assign n4830 = n2777 ? encrypted_data_buf[726] : n4822;   // modexp_top.v(481)
    assign n4831 = n2777 ? encrypted_data_buf[725] : n4823;   // modexp_top.v(481)
    assign n4832 = n2777 ? encrypted_data_buf[724] : n4824;   // modexp_top.v(481)
    assign n4833 = n2777 ? encrypted_data_buf[723] : n4825;   // modexp_top.v(481)
    assign n4834 = n2777 ? encrypted_data_buf[722] : n4826;   // modexp_top.v(481)
    assign n4835 = n2777 ? encrypted_data_buf[721] : n4827;   // modexp_top.v(481)
    assign n4836 = n2777 ? encrypted_data_buf[720] : n4828;   // modexp_top.v(481)
    assign n4837 = n2772 ? encrypted_data_buf[719] : n4829;   // modexp_top.v(481)
    assign n4838 = n2772 ? encrypted_data_buf[718] : n4830;   // modexp_top.v(481)
    assign n4839 = n2772 ? encrypted_data_buf[717] : n4831;   // modexp_top.v(481)
    assign n4840 = n2772 ? encrypted_data_buf[716] : n4832;   // modexp_top.v(481)
    assign n4841 = n2772 ? encrypted_data_buf[715] : n4833;   // modexp_top.v(481)
    assign n4842 = n2772 ? encrypted_data_buf[714] : n4834;   // modexp_top.v(481)
    assign n4843 = n2772 ? encrypted_data_buf[713] : n4835;   // modexp_top.v(481)
    assign n4844 = n2772 ? encrypted_data_buf[712] : n4836;   // modexp_top.v(481)
    assign n4845 = n2767 ? encrypted_data_buf[711] : n4837;   // modexp_top.v(481)
    assign n4846 = n2767 ? encrypted_data_buf[710] : n4838;   // modexp_top.v(481)
    assign n4847 = n2767 ? encrypted_data_buf[709] : n4839;   // modexp_top.v(481)
    assign n4848 = n2767 ? encrypted_data_buf[708] : n4840;   // modexp_top.v(481)
    assign n4849 = n2767 ? encrypted_data_buf[707] : n4841;   // modexp_top.v(481)
    assign n4850 = n2767 ? encrypted_data_buf[706] : n4842;   // modexp_top.v(481)
    assign n4851 = n2767 ? encrypted_data_buf[705] : n4843;   // modexp_top.v(481)
    assign n4852 = n2767 ? encrypted_data_buf[704] : n4844;   // modexp_top.v(481)
    assign n4853 = n2761 ? encrypted_data_buf[703] : n4845;   // modexp_top.v(481)
    assign n4854 = n2761 ? encrypted_data_buf[702] : n4846;   // modexp_top.v(481)
    assign n4855 = n2761 ? encrypted_data_buf[701] : n4847;   // modexp_top.v(481)
    assign n4856 = n2761 ? encrypted_data_buf[700] : n4848;   // modexp_top.v(481)
    assign n4857 = n2761 ? encrypted_data_buf[699] : n4849;   // modexp_top.v(481)
    assign n4858 = n2761 ? encrypted_data_buf[698] : n4850;   // modexp_top.v(481)
    assign n4859 = n2761 ? encrypted_data_buf[697] : n4851;   // modexp_top.v(481)
    assign n4860 = n2761 ? encrypted_data_buf[696] : n4852;   // modexp_top.v(481)
    assign n4861 = n2757 ? encrypted_data_buf[695] : n4853;   // modexp_top.v(481)
    assign n4862 = n2757 ? encrypted_data_buf[694] : n4854;   // modexp_top.v(481)
    assign n4863 = n2757 ? encrypted_data_buf[693] : n4855;   // modexp_top.v(481)
    assign n4864 = n2757 ? encrypted_data_buf[692] : n4856;   // modexp_top.v(481)
    assign n4865 = n2757 ? encrypted_data_buf[691] : n4857;   // modexp_top.v(481)
    assign n4866 = n2757 ? encrypted_data_buf[690] : n4858;   // modexp_top.v(481)
    assign n4867 = n2757 ? encrypted_data_buf[689] : n4859;   // modexp_top.v(481)
    assign n4868 = n2757 ? encrypted_data_buf[688] : n4860;   // modexp_top.v(481)
    assign n4869 = n2752 ? encrypted_data_buf[687] : n4861;   // modexp_top.v(481)
    assign n4870 = n2752 ? encrypted_data_buf[686] : n4862;   // modexp_top.v(481)
    assign n4871 = n2752 ? encrypted_data_buf[685] : n4863;   // modexp_top.v(481)
    assign n4872 = n2752 ? encrypted_data_buf[684] : n4864;   // modexp_top.v(481)
    assign n4873 = n2752 ? encrypted_data_buf[683] : n4865;   // modexp_top.v(481)
    assign n4874 = n2752 ? encrypted_data_buf[682] : n4866;   // modexp_top.v(481)
    assign n4875 = n2752 ? encrypted_data_buf[681] : n4867;   // modexp_top.v(481)
    assign n4876 = n2752 ? encrypted_data_buf[680] : n4868;   // modexp_top.v(481)
    assign n4877 = n2747 ? encrypted_data_buf[679] : n4869;   // modexp_top.v(481)
    assign n4878 = n2747 ? encrypted_data_buf[678] : n4870;   // modexp_top.v(481)
    assign n4879 = n2747 ? encrypted_data_buf[677] : n4871;   // modexp_top.v(481)
    assign n4880 = n2747 ? encrypted_data_buf[676] : n4872;   // modexp_top.v(481)
    assign n4881 = n2747 ? encrypted_data_buf[675] : n4873;   // modexp_top.v(481)
    assign n4882 = n2747 ? encrypted_data_buf[674] : n4874;   // modexp_top.v(481)
    assign n4883 = n2747 ? encrypted_data_buf[673] : n4875;   // modexp_top.v(481)
    assign n4884 = n2747 ? encrypted_data_buf[672] : n4876;   // modexp_top.v(481)
    assign n4885 = n2741 ? encrypted_data_buf[671] : n4877;   // modexp_top.v(481)
    assign n4886 = n2741 ? encrypted_data_buf[670] : n4878;   // modexp_top.v(481)
    assign n4887 = n2741 ? encrypted_data_buf[669] : n4879;   // modexp_top.v(481)
    assign n4888 = n2741 ? encrypted_data_buf[668] : n4880;   // modexp_top.v(481)
    assign n4889 = n2741 ? encrypted_data_buf[667] : n4881;   // modexp_top.v(481)
    assign n4890 = n2741 ? encrypted_data_buf[666] : n4882;   // modexp_top.v(481)
    assign n4891 = n2741 ? encrypted_data_buf[665] : n4883;   // modexp_top.v(481)
    assign n4892 = n2741 ? encrypted_data_buf[664] : n4884;   // modexp_top.v(481)
    assign n4893 = n2736 ? encrypted_data_buf[663] : n4885;   // modexp_top.v(481)
    assign n4894 = n2736 ? encrypted_data_buf[662] : n4886;   // modexp_top.v(481)
    assign n4895 = n2736 ? encrypted_data_buf[661] : n4887;   // modexp_top.v(481)
    assign n4896 = n2736 ? encrypted_data_buf[660] : n4888;   // modexp_top.v(481)
    assign n4897 = n2736 ? encrypted_data_buf[659] : n4889;   // modexp_top.v(481)
    assign n4898 = n2736 ? encrypted_data_buf[658] : n4890;   // modexp_top.v(481)
    assign n4899 = n2736 ? encrypted_data_buf[657] : n4891;   // modexp_top.v(481)
    assign n4900 = n2736 ? encrypted_data_buf[656] : n4892;   // modexp_top.v(481)
    assign n4901 = n2730 ? encrypted_data_buf[655] : n4893;   // modexp_top.v(481)
    assign n4902 = n2730 ? encrypted_data_buf[654] : n4894;   // modexp_top.v(481)
    assign n4903 = n2730 ? encrypted_data_buf[653] : n4895;   // modexp_top.v(481)
    assign n4904 = n2730 ? encrypted_data_buf[652] : n4896;   // modexp_top.v(481)
    assign n4905 = n2730 ? encrypted_data_buf[651] : n4897;   // modexp_top.v(481)
    assign n4906 = n2730 ? encrypted_data_buf[650] : n4898;   // modexp_top.v(481)
    assign n4907 = n2730 ? encrypted_data_buf[649] : n4899;   // modexp_top.v(481)
    assign n4908 = n2730 ? encrypted_data_buf[648] : n4900;   // modexp_top.v(481)
    assign n4909 = n2724 ? encrypted_data_buf[647] : n4901;   // modexp_top.v(481)
    assign n4910 = n2724 ? encrypted_data_buf[646] : n4902;   // modexp_top.v(481)
    assign n4911 = n2724 ? encrypted_data_buf[645] : n4903;   // modexp_top.v(481)
    assign n4912 = n2724 ? encrypted_data_buf[644] : n4904;   // modexp_top.v(481)
    assign n4913 = n2724 ? encrypted_data_buf[643] : n4905;   // modexp_top.v(481)
    assign n4914 = n2724 ? encrypted_data_buf[642] : n4906;   // modexp_top.v(481)
    assign n4915 = n2724 ? encrypted_data_buf[641] : n4907;   // modexp_top.v(481)
    assign n4916 = n2724 ? encrypted_data_buf[640] : n4908;   // modexp_top.v(481)
    assign n4917 = n2717 ? encrypted_data_buf[639] : n4909;   // modexp_top.v(481)
    assign n4918 = n2717 ? encrypted_data_buf[638] : n4910;   // modexp_top.v(481)
    assign n4919 = n2717 ? encrypted_data_buf[637] : n4911;   // modexp_top.v(481)
    assign n4920 = n2717 ? encrypted_data_buf[636] : n4912;   // modexp_top.v(481)
    assign n4921 = n2717 ? encrypted_data_buf[635] : n4913;   // modexp_top.v(481)
    assign n4922 = n2717 ? encrypted_data_buf[634] : n4914;   // modexp_top.v(481)
    assign n4923 = n2717 ? encrypted_data_buf[633] : n4915;   // modexp_top.v(481)
    assign n4924 = n2717 ? encrypted_data_buf[632] : n4916;   // modexp_top.v(481)
    assign n4925 = n2713 ? encrypted_data_buf[631] : n4917;   // modexp_top.v(481)
    assign n4926 = n2713 ? encrypted_data_buf[630] : n4918;   // modexp_top.v(481)
    assign n4927 = n2713 ? encrypted_data_buf[629] : n4919;   // modexp_top.v(481)
    assign n4928 = n2713 ? encrypted_data_buf[628] : n4920;   // modexp_top.v(481)
    assign n4929 = n2713 ? encrypted_data_buf[627] : n4921;   // modexp_top.v(481)
    assign n4930 = n2713 ? encrypted_data_buf[626] : n4922;   // modexp_top.v(481)
    assign n4931 = n2713 ? encrypted_data_buf[625] : n4923;   // modexp_top.v(481)
    assign n4932 = n2713 ? encrypted_data_buf[624] : n4924;   // modexp_top.v(481)
    assign n4933 = n2708 ? encrypted_data_buf[623] : n4925;   // modexp_top.v(481)
    assign n4934 = n2708 ? encrypted_data_buf[622] : n4926;   // modexp_top.v(481)
    assign n4935 = n2708 ? encrypted_data_buf[621] : n4927;   // modexp_top.v(481)
    assign n4936 = n2708 ? encrypted_data_buf[620] : n4928;   // modexp_top.v(481)
    assign n4937 = n2708 ? encrypted_data_buf[619] : n4929;   // modexp_top.v(481)
    assign n4938 = n2708 ? encrypted_data_buf[618] : n4930;   // modexp_top.v(481)
    assign n4939 = n2708 ? encrypted_data_buf[617] : n4931;   // modexp_top.v(481)
    assign n4940 = n2708 ? encrypted_data_buf[616] : n4932;   // modexp_top.v(481)
    assign n4941 = n2703 ? encrypted_data_buf[615] : n4933;   // modexp_top.v(481)
    assign n4942 = n2703 ? encrypted_data_buf[614] : n4934;   // modexp_top.v(481)
    assign n4943 = n2703 ? encrypted_data_buf[613] : n4935;   // modexp_top.v(481)
    assign n4944 = n2703 ? encrypted_data_buf[612] : n4936;   // modexp_top.v(481)
    assign n4945 = n2703 ? encrypted_data_buf[611] : n4937;   // modexp_top.v(481)
    assign n4946 = n2703 ? encrypted_data_buf[610] : n4938;   // modexp_top.v(481)
    assign n4947 = n2703 ? encrypted_data_buf[609] : n4939;   // modexp_top.v(481)
    assign n4948 = n2703 ? encrypted_data_buf[608] : n4940;   // modexp_top.v(481)
    assign n4949 = n2697 ? encrypted_data_buf[607] : n4941;   // modexp_top.v(481)
    assign n4950 = n2697 ? encrypted_data_buf[606] : n4942;   // modexp_top.v(481)
    assign n4951 = n2697 ? encrypted_data_buf[605] : n4943;   // modexp_top.v(481)
    assign n4952 = n2697 ? encrypted_data_buf[604] : n4944;   // modexp_top.v(481)
    assign n4953 = n2697 ? encrypted_data_buf[603] : n4945;   // modexp_top.v(481)
    assign n4954 = n2697 ? encrypted_data_buf[602] : n4946;   // modexp_top.v(481)
    assign n4955 = n2697 ? encrypted_data_buf[601] : n4947;   // modexp_top.v(481)
    assign n4956 = n2697 ? encrypted_data_buf[600] : n4948;   // modexp_top.v(481)
    assign n4957 = n2692 ? encrypted_data_buf[599] : n4949;   // modexp_top.v(481)
    assign n4958 = n2692 ? encrypted_data_buf[598] : n4950;   // modexp_top.v(481)
    assign n4959 = n2692 ? encrypted_data_buf[597] : n4951;   // modexp_top.v(481)
    assign n4960 = n2692 ? encrypted_data_buf[596] : n4952;   // modexp_top.v(481)
    assign n4961 = n2692 ? encrypted_data_buf[595] : n4953;   // modexp_top.v(481)
    assign n4962 = n2692 ? encrypted_data_buf[594] : n4954;   // modexp_top.v(481)
    assign n4963 = n2692 ? encrypted_data_buf[593] : n4955;   // modexp_top.v(481)
    assign n4964 = n2692 ? encrypted_data_buf[592] : n4956;   // modexp_top.v(481)
    assign n4965 = n2686 ? encrypted_data_buf[591] : n4957;   // modexp_top.v(481)
    assign n4966 = n2686 ? encrypted_data_buf[590] : n4958;   // modexp_top.v(481)
    assign n4967 = n2686 ? encrypted_data_buf[589] : n4959;   // modexp_top.v(481)
    assign n4968 = n2686 ? encrypted_data_buf[588] : n4960;   // modexp_top.v(481)
    assign n4969 = n2686 ? encrypted_data_buf[587] : n4961;   // modexp_top.v(481)
    assign n4970 = n2686 ? encrypted_data_buf[586] : n4962;   // modexp_top.v(481)
    assign n4971 = n2686 ? encrypted_data_buf[585] : n4963;   // modexp_top.v(481)
    assign n4972 = n2686 ? encrypted_data_buf[584] : n4964;   // modexp_top.v(481)
    assign n4973 = n2680 ? encrypted_data_buf[583] : n4965;   // modexp_top.v(481)
    assign n4974 = n2680 ? encrypted_data_buf[582] : n4966;   // modexp_top.v(481)
    assign n4975 = n2680 ? encrypted_data_buf[581] : n4967;   // modexp_top.v(481)
    assign n4976 = n2680 ? encrypted_data_buf[580] : n4968;   // modexp_top.v(481)
    assign n4977 = n2680 ? encrypted_data_buf[579] : n4969;   // modexp_top.v(481)
    assign n4978 = n2680 ? encrypted_data_buf[578] : n4970;   // modexp_top.v(481)
    assign n4979 = n2680 ? encrypted_data_buf[577] : n4971;   // modexp_top.v(481)
    assign n4980 = n2680 ? encrypted_data_buf[576] : n4972;   // modexp_top.v(481)
    assign n4981 = n2673 ? encrypted_data_buf[575] : n4973;   // modexp_top.v(481)
    assign n4982 = n2673 ? encrypted_data_buf[574] : n4974;   // modexp_top.v(481)
    assign n4983 = n2673 ? encrypted_data_buf[573] : n4975;   // modexp_top.v(481)
    assign n4984 = n2673 ? encrypted_data_buf[572] : n4976;   // modexp_top.v(481)
    assign n4985 = n2673 ? encrypted_data_buf[571] : n4977;   // modexp_top.v(481)
    assign n4986 = n2673 ? encrypted_data_buf[570] : n4978;   // modexp_top.v(481)
    assign n4987 = n2673 ? encrypted_data_buf[569] : n4979;   // modexp_top.v(481)
    assign n4988 = n2673 ? encrypted_data_buf[568] : n4980;   // modexp_top.v(481)
    assign n4989 = n2668 ? encrypted_data_buf[567] : n4981;   // modexp_top.v(481)
    assign n4990 = n2668 ? encrypted_data_buf[566] : n4982;   // modexp_top.v(481)
    assign n4991 = n2668 ? encrypted_data_buf[565] : n4983;   // modexp_top.v(481)
    assign n4992 = n2668 ? encrypted_data_buf[564] : n4984;   // modexp_top.v(481)
    assign n4993 = n2668 ? encrypted_data_buf[563] : n4985;   // modexp_top.v(481)
    assign n4994 = n2668 ? encrypted_data_buf[562] : n4986;   // modexp_top.v(481)
    assign n4995 = n2668 ? encrypted_data_buf[561] : n4987;   // modexp_top.v(481)
    assign n4996 = n2668 ? encrypted_data_buf[560] : n4988;   // modexp_top.v(481)
    assign n4997 = n2662 ? encrypted_data_buf[559] : n4989;   // modexp_top.v(481)
    assign n4998 = n2662 ? encrypted_data_buf[558] : n4990;   // modexp_top.v(481)
    assign n4999 = n2662 ? encrypted_data_buf[557] : n4991;   // modexp_top.v(481)
    assign n5000 = n2662 ? encrypted_data_buf[556] : n4992;   // modexp_top.v(481)
    assign n5001 = n2662 ? encrypted_data_buf[555] : n4993;   // modexp_top.v(481)
    assign n5002 = n2662 ? encrypted_data_buf[554] : n4994;   // modexp_top.v(481)
    assign n5003 = n2662 ? encrypted_data_buf[553] : n4995;   // modexp_top.v(481)
    assign n5004 = n2662 ? encrypted_data_buf[552] : n4996;   // modexp_top.v(481)
    assign n5005 = n2656 ? encrypted_data_buf[551] : n4997;   // modexp_top.v(481)
    assign n5006 = n2656 ? encrypted_data_buf[550] : n4998;   // modexp_top.v(481)
    assign n5007 = n2656 ? encrypted_data_buf[549] : n4999;   // modexp_top.v(481)
    assign n5008 = n2656 ? encrypted_data_buf[548] : n5000;   // modexp_top.v(481)
    assign n5009 = n2656 ? encrypted_data_buf[547] : n5001;   // modexp_top.v(481)
    assign n5010 = n2656 ? encrypted_data_buf[546] : n5002;   // modexp_top.v(481)
    assign n5011 = n2656 ? encrypted_data_buf[545] : n5003;   // modexp_top.v(481)
    assign n5012 = n2656 ? encrypted_data_buf[544] : n5004;   // modexp_top.v(481)
    assign n5013 = n2649 ? encrypted_data_buf[543] : n5005;   // modexp_top.v(481)
    assign n5014 = n2649 ? encrypted_data_buf[542] : n5006;   // modexp_top.v(481)
    assign n5015 = n2649 ? encrypted_data_buf[541] : n5007;   // modexp_top.v(481)
    assign n5016 = n2649 ? encrypted_data_buf[540] : n5008;   // modexp_top.v(481)
    assign n5017 = n2649 ? encrypted_data_buf[539] : n5009;   // modexp_top.v(481)
    assign n5018 = n2649 ? encrypted_data_buf[538] : n5010;   // modexp_top.v(481)
    assign n5019 = n2649 ? encrypted_data_buf[537] : n5011;   // modexp_top.v(481)
    assign n5020 = n2649 ? encrypted_data_buf[536] : n5012;   // modexp_top.v(481)
    assign n5021 = n2643 ? encrypted_data_buf[535] : n5013;   // modexp_top.v(481)
    assign n5022 = n2643 ? encrypted_data_buf[534] : n5014;   // modexp_top.v(481)
    assign n5023 = n2643 ? encrypted_data_buf[533] : n5015;   // modexp_top.v(481)
    assign n5024 = n2643 ? encrypted_data_buf[532] : n5016;   // modexp_top.v(481)
    assign n5025 = n2643 ? encrypted_data_buf[531] : n5017;   // modexp_top.v(481)
    assign n5026 = n2643 ? encrypted_data_buf[530] : n5018;   // modexp_top.v(481)
    assign n5027 = n2643 ? encrypted_data_buf[529] : n5019;   // modexp_top.v(481)
    assign n5028 = n2643 ? encrypted_data_buf[528] : n5020;   // modexp_top.v(481)
    assign n5029 = n2636 ? encrypted_data_buf[527] : n5021;   // modexp_top.v(481)
    assign n5030 = n2636 ? encrypted_data_buf[526] : n5022;   // modexp_top.v(481)
    assign n5031 = n2636 ? encrypted_data_buf[525] : n5023;   // modexp_top.v(481)
    assign n5032 = n2636 ? encrypted_data_buf[524] : n5024;   // modexp_top.v(481)
    assign n5033 = n2636 ? encrypted_data_buf[523] : n5025;   // modexp_top.v(481)
    assign n5034 = n2636 ? encrypted_data_buf[522] : n5026;   // modexp_top.v(481)
    assign n5035 = n2636 ? encrypted_data_buf[521] : n5027;   // modexp_top.v(481)
    assign n5036 = n2636 ? encrypted_data_buf[520] : n5028;   // modexp_top.v(481)
    assign n5037 = n2629 ? encrypted_data_buf[519] : n5029;   // modexp_top.v(481)
    assign n5038 = n2629 ? encrypted_data_buf[518] : n5030;   // modexp_top.v(481)
    assign n5039 = n2629 ? encrypted_data_buf[517] : n5031;   // modexp_top.v(481)
    assign n5040 = n2629 ? encrypted_data_buf[516] : n5032;   // modexp_top.v(481)
    assign n5041 = n2629 ? encrypted_data_buf[515] : n5033;   // modexp_top.v(481)
    assign n5042 = n2629 ? encrypted_data_buf[514] : n5034;   // modexp_top.v(481)
    assign n5043 = n2629 ? encrypted_data_buf[513] : n5035;   // modexp_top.v(481)
    assign n5044 = n2629 ? encrypted_data_buf[512] : n5036;   // modexp_top.v(481)
    assign n5045 = n2621 ? encrypted_data_buf[511] : n5037;   // modexp_top.v(481)
    assign n5046 = n2621 ? encrypted_data_buf[510] : n5038;   // modexp_top.v(481)
    assign n5047 = n2621 ? encrypted_data_buf[509] : n5039;   // modexp_top.v(481)
    assign n5048 = n2621 ? encrypted_data_buf[508] : n5040;   // modexp_top.v(481)
    assign n5049 = n2621 ? encrypted_data_buf[507] : n5041;   // modexp_top.v(481)
    assign n5050 = n2621 ? encrypted_data_buf[506] : n5042;   // modexp_top.v(481)
    assign n5051 = n2621 ? encrypted_data_buf[505] : n5043;   // modexp_top.v(481)
    assign n5052 = n2621 ? encrypted_data_buf[504] : n5044;   // modexp_top.v(481)
    assign n5053 = n2618 ? encrypted_data_buf[503] : n5045;   // modexp_top.v(481)
    assign n5054 = n2618 ? encrypted_data_buf[502] : n5046;   // modexp_top.v(481)
    assign n5055 = n2618 ? encrypted_data_buf[501] : n5047;   // modexp_top.v(481)
    assign n5056 = n2618 ? encrypted_data_buf[500] : n5048;   // modexp_top.v(481)
    assign n5057 = n2618 ? encrypted_data_buf[499] : n5049;   // modexp_top.v(481)
    assign n5058 = n2618 ? encrypted_data_buf[498] : n5050;   // modexp_top.v(481)
    assign n5059 = n2618 ? encrypted_data_buf[497] : n5051;   // modexp_top.v(481)
    assign n5060 = n2618 ? encrypted_data_buf[496] : n5052;   // modexp_top.v(481)
    assign n5061 = n2614 ? encrypted_data_buf[495] : n5053;   // modexp_top.v(481)
    assign n5062 = n2614 ? encrypted_data_buf[494] : n5054;   // modexp_top.v(481)
    assign n5063 = n2614 ? encrypted_data_buf[493] : n5055;   // modexp_top.v(481)
    assign n5064 = n2614 ? encrypted_data_buf[492] : n5056;   // modexp_top.v(481)
    assign n5065 = n2614 ? encrypted_data_buf[491] : n5057;   // modexp_top.v(481)
    assign n5066 = n2614 ? encrypted_data_buf[490] : n5058;   // modexp_top.v(481)
    assign n5067 = n2614 ? encrypted_data_buf[489] : n5059;   // modexp_top.v(481)
    assign n5068 = n2614 ? encrypted_data_buf[488] : n5060;   // modexp_top.v(481)
    assign n5069 = n2610 ? encrypted_data_buf[487] : n5061;   // modexp_top.v(481)
    assign n5070 = n2610 ? encrypted_data_buf[486] : n5062;   // modexp_top.v(481)
    assign n5071 = n2610 ? encrypted_data_buf[485] : n5063;   // modexp_top.v(481)
    assign n5072 = n2610 ? encrypted_data_buf[484] : n5064;   // modexp_top.v(481)
    assign n5073 = n2610 ? encrypted_data_buf[483] : n5065;   // modexp_top.v(481)
    assign n5074 = n2610 ? encrypted_data_buf[482] : n5066;   // modexp_top.v(481)
    assign n5075 = n2610 ? encrypted_data_buf[481] : n5067;   // modexp_top.v(481)
    assign n5076 = n2610 ? encrypted_data_buf[480] : n5068;   // modexp_top.v(481)
    assign n5077 = n2605 ? encrypted_data_buf[479] : n5069;   // modexp_top.v(481)
    assign n5078 = n2605 ? encrypted_data_buf[478] : n5070;   // modexp_top.v(481)
    assign n5079 = n2605 ? encrypted_data_buf[477] : n5071;   // modexp_top.v(481)
    assign n5080 = n2605 ? encrypted_data_buf[476] : n5072;   // modexp_top.v(481)
    assign n5081 = n2605 ? encrypted_data_buf[475] : n5073;   // modexp_top.v(481)
    assign n5082 = n2605 ? encrypted_data_buf[474] : n5074;   // modexp_top.v(481)
    assign n5083 = n2605 ? encrypted_data_buf[473] : n5075;   // modexp_top.v(481)
    assign n5084 = n2605 ? encrypted_data_buf[472] : n5076;   // modexp_top.v(481)
    assign n5085 = n2601 ? encrypted_data_buf[471] : n5077;   // modexp_top.v(481)
    assign n5086 = n2601 ? encrypted_data_buf[470] : n5078;   // modexp_top.v(481)
    assign n5087 = n2601 ? encrypted_data_buf[469] : n5079;   // modexp_top.v(481)
    assign n5088 = n2601 ? encrypted_data_buf[468] : n5080;   // modexp_top.v(481)
    assign n5089 = n2601 ? encrypted_data_buf[467] : n5081;   // modexp_top.v(481)
    assign n5090 = n2601 ? encrypted_data_buf[466] : n5082;   // modexp_top.v(481)
    assign n5091 = n2601 ? encrypted_data_buf[465] : n5083;   // modexp_top.v(481)
    assign n5092 = n2601 ? encrypted_data_buf[464] : n5084;   // modexp_top.v(481)
    assign n5093 = n2596 ? encrypted_data_buf[463] : n5085;   // modexp_top.v(481)
    assign n5094 = n2596 ? encrypted_data_buf[462] : n5086;   // modexp_top.v(481)
    assign n5095 = n2596 ? encrypted_data_buf[461] : n5087;   // modexp_top.v(481)
    assign n5096 = n2596 ? encrypted_data_buf[460] : n5088;   // modexp_top.v(481)
    assign n5097 = n2596 ? encrypted_data_buf[459] : n5089;   // modexp_top.v(481)
    assign n5098 = n2596 ? encrypted_data_buf[458] : n5090;   // modexp_top.v(481)
    assign n5099 = n2596 ? encrypted_data_buf[457] : n5091;   // modexp_top.v(481)
    assign n5100 = n2596 ? encrypted_data_buf[456] : n5092;   // modexp_top.v(481)
    assign n5101 = n2591 ? encrypted_data_buf[455] : n5093;   // modexp_top.v(481)
    assign n5102 = n2591 ? encrypted_data_buf[454] : n5094;   // modexp_top.v(481)
    assign n5103 = n2591 ? encrypted_data_buf[453] : n5095;   // modexp_top.v(481)
    assign n5104 = n2591 ? encrypted_data_buf[452] : n5096;   // modexp_top.v(481)
    assign n5105 = n2591 ? encrypted_data_buf[451] : n5097;   // modexp_top.v(481)
    assign n5106 = n2591 ? encrypted_data_buf[450] : n5098;   // modexp_top.v(481)
    assign n5107 = n2591 ? encrypted_data_buf[449] : n5099;   // modexp_top.v(481)
    assign n5108 = n2591 ? encrypted_data_buf[448] : n5100;   // modexp_top.v(481)
    assign n5109 = n2585 ? encrypted_data_buf[447] : n5101;   // modexp_top.v(481)
    assign n5110 = n2585 ? encrypted_data_buf[446] : n5102;   // modexp_top.v(481)
    assign n5111 = n2585 ? encrypted_data_buf[445] : n5103;   // modexp_top.v(481)
    assign n5112 = n2585 ? encrypted_data_buf[444] : n5104;   // modexp_top.v(481)
    assign n5113 = n2585 ? encrypted_data_buf[443] : n5105;   // modexp_top.v(481)
    assign n5114 = n2585 ? encrypted_data_buf[442] : n5106;   // modexp_top.v(481)
    assign n5115 = n2585 ? encrypted_data_buf[441] : n5107;   // modexp_top.v(481)
    assign n5116 = n2585 ? encrypted_data_buf[440] : n5108;   // modexp_top.v(481)
    assign n5117 = n2581 ? encrypted_data_buf[439] : n5109;   // modexp_top.v(481)
    assign n5118 = n2581 ? encrypted_data_buf[438] : n5110;   // modexp_top.v(481)
    assign n5119 = n2581 ? encrypted_data_buf[437] : n5111;   // modexp_top.v(481)
    assign n5120 = n2581 ? encrypted_data_buf[436] : n5112;   // modexp_top.v(481)
    assign n5121 = n2581 ? encrypted_data_buf[435] : n5113;   // modexp_top.v(481)
    assign n5122 = n2581 ? encrypted_data_buf[434] : n5114;   // modexp_top.v(481)
    assign n5123 = n2581 ? encrypted_data_buf[433] : n5115;   // modexp_top.v(481)
    assign n5124 = n2581 ? encrypted_data_buf[432] : n5116;   // modexp_top.v(481)
    assign n5125 = n2576 ? encrypted_data_buf[431] : n5117;   // modexp_top.v(481)
    assign n5126 = n2576 ? encrypted_data_buf[430] : n5118;   // modexp_top.v(481)
    assign n5127 = n2576 ? encrypted_data_buf[429] : n5119;   // modexp_top.v(481)
    assign n5128 = n2576 ? encrypted_data_buf[428] : n5120;   // modexp_top.v(481)
    assign n5129 = n2576 ? encrypted_data_buf[427] : n5121;   // modexp_top.v(481)
    assign n5130 = n2576 ? encrypted_data_buf[426] : n5122;   // modexp_top.v(481)
    assign n5131 = n2576 ? encrypted_data_buf[425] : n5123;   // modexp_top.v(481)
    assign n5132 = n2576 ? encrypted_data_buf[424] : n5124;   // modexp_top.v(481)
    assign n5133 = n2571 ? encrypted_data_buf[423] : n5125;   // modexp_top.v(481)
    assign n5134 = n2571 ? encrypted_data_buf[422] : n5126;   // modexp_top.v(481)
    assign n5135 = n2571 ? encrypted_data_buf[421] : n5127;   // modexp_top.v(481)
    assign n5136 = n2571 ? encrypted_data_buf[420] : n5128;   // modexp_top.v(481)
    assign n5137 = n2571 ? encrypted_data_buf[419] : n5129;   // modexp_top.v(481)
    assign n5138 = n2571 ? encrypted_data_buf[418] : n5130;   // modexp_top.v(481)
    assign n5139 = n2571 ? encrypted_data_buf[417] : n5131;   // modexp_top.v(481)
    assign n5140 = n2571 ? encrypted_data_buf[416] : n5132;   // modexp_top.v(481)
    assign n5141 = n2565 ? encrypted_data_buf[415] : n5133;   // modexp_top.v(481)
    assign n5142 = n2565 ? encrypted_data_buf[414] : n5134;   // modexp_top.v(481)
    assign n5143 = n2565 ? encrypted_data_buf[413] : n5135;   // modexp_top.v(481)
    assign n5144 = n2565 ? encrypted_data_buf[412] : n5136;   // modexp_top.v(481)
    assign n5145 = n2565 ? encrypted_data_buf[411] : n5137;   // modexp_top.v(481)
    assign n5146 = n2565 ? encrypted_data_buf[410] : n5138;   // modexp_top.v(481)
    assign n5147 = n2565 ? encrypted_data_buf[409] : n5139;   // modexp_top.v(481)
    assign n5148 = n2565 ? encrypted_data_buf[408] : n5140;   // modexp_top.v(481)
    assign n5149 = n2560 ? encrypted_data_buf[407] : n5141;   // modexp_top.v(481)
    assign n5150 = n2560 ? encrypted_data_buf[406] : n5142;   // modexp_top.v(481)
    assign n5151 = n2560 ? encrypted_data_buf[405] : n5143;   // modexp_top.v(481)
    assign n5152 = n2560 ? encrypted_data_buf[404] : n5144;   // modexp_top.v(481)
    assign n5153 = n2560 ? encrypted_data_buf[403] : n5145;   // modexp_top.v(481)
    assign n5154 = n2560 ? encrypted_data_buf[402] : n5146;   // modexp_top.v(481)
    assign n5155 = n2560 ? encrypted_data_buf[401] : n5147;   // modexp_top.v(481)
    assign n5156 = n2560 ? encrypted_data_buf[400] : n5148;   // modexp_top.v(481)
    assign n5157 = n2554 ? encrypted_data_buf[399] : n5149;   // modexp_top.v(481)
    assign n5158 = n2554 ? encrypted_data_buf[398] : n5150;   // modexp_top.v(481)
    assign n5159 = n2554 ? encrypted_data_buf[397] : n5151;   // modexp_top.v(481)
    assign n5160 = n2554 ? encrypted_data_buf[396] : n5152;   // modexp_top.v(481)
    assign n5161 = n2554 ? encrypted_data_buf[395] : n5153;   // modexp_top.v(481)
    assign n5162 = n2554 ? encrypted_data_buf[394] : n5154;   // modexp_top.v(481)
    assign n5163 = n2554 ? encrypted_data_buf[393] : n5155;   // modexp_top.v(481)
    assign n5164 = n2554 ? encrypted_data_buf[392] : n5156;   // modexp_top.v(481)
    assign n5165 = n2548 ? encrypted_data_buf[391] : n5157;   // modexp_top.v(481)
    assign n5166 = n2548 ? encrypted_data_buf[390] : n5158;   // modexp_top.v(481)
    assign n5167 = n2548 ? encrypted_data_buf[389] : n5159;   // modexp_top.v(481)
    assign n5168 = n2548 ? encrypted_data_buf[388] : n5160;   // modexp_top.v(481)
    assign n5169 = n2548 ? encrypted_data_buf[387] : n5161;   // modexp_top.v(481)
    assign n5170 = n2548 ? encrypted_data_buf[386] : n5162;   // modexp_top.v(481)
    assign n5171 = n2548 ? encrypted_data_buf[385] : n5163;   // modexp_top.v(481)
    assign n5172 = n2548 ? encrypted_data_buf[384] : n5164;   // modexp_top.v(481)
    assign n5173 = n2541 ? encrypted_data_buf[383] : n5165;   // modexp_top.v(481)
    assign n5174 = n2541 ? encrypted_data_buf[382] : n5166;   // modexp_top.v(481)
    assign n5175 = n2541 ? encrypted_data_buf[381] : n5167;   // modexp_top.v(481)
    assign n5176 = n2541 ? encrypted_data_buf[380] : n5168;   // modexp_top.v(481)
    assign n5177 = n2541 ? encrypted_data_buf[379] : n5169;   // modexp_top.v(481)
    assign n5178 = n2541 ? encrypted_data_buf[378] : n5170;   // modexp_top.v(481)
    assign n5179 = n2541 ? encrypted_data_buf[377] : n5171;   // modexp_top.v(481)
    assign n5180 = n2541 ? encrypted_data_buf[376] : n5172;   // modexp_top.v(481)
    assign n5181 = n2537 ? encrypted_data_buf[375] : n5173;   // modexp_top.v(481)
    assign n5182 = n2537 ? encrypted_data_buf[374] : n5174;   // modexp_top.v(481)
    assign n5183 = n2537 ? encrypted_data_buf[373] : n5175;   // modexp_top.v(481)
    assign n5184 = n2537 ? encrypted_data_buf[372] : n5176;   // modexp_top.v(481)
    assign n5185 = n2537 ? encrypted_data_buf[371] : n5177;   // modexp_top.v(481)
    assign n5186 = n2537 ? encrypted_data_buf[370] : n5178;   // modexp_top.v(481)
    assign n5187 = n2537 ? encrypted_data_buf[369] : n5179;   // modexp_top.v(481)
    assign n5188 = n2537 ? encrypted_data_buf[368] : n5180;   // modexp_top.v(481)
    assign n5189 = n2532 ? encrypted_data_buf[367] : n5181;   // modexp_top.v(481)
    assign n5190 = n2532 ? encrypted_data_buf[366] : n5182;   // modexp_top.v(481)
    assign n5191 = n2532 ? encrypted_data_buf[365] : n5183;   // modexp_top.v(481)
    assign n5192 = n2532 ? encrypted_data_buf[364] : n5184;   // modexp_top.v(481)
    assign n5193 = n2532 ? encrypted_data_buf[363] : n5185;   // modexp_top.v(481)
    assign n5194 = n2532 ? encrypted_data_buf[362] : n5186;   // modexp_top.v(481)
    assign n5195 = n2532 ? encrypted_data_buf[361] : n5187;   // modexp_top.v(481)
    assign n5196 = n2532 ? encrypted_data_buf[360] : n5188;   // modexp_top.v(481)
    assign n5197 = n2527 ? encrypted_data_buf[359] : n5189;   // modexp_top.v(481)
    assign n5198 = n2527 ? encrypted_data_buf[358] : n5190;   // modexp_top.v(481)
    assign n5199 = n2527 ? encrypted_data_buf[357] : n5191;   // modexp_top.v(481)
    assign n5200 = n2527 ? encrypted_data_buf[356] : n5192;   // modexp_top.v(481)
    assign n5201 = n2527 ? encrypted_data_buf[355] : n5193;   // modexp_top.v(481)
    assign n5202 = n2527 ? encrypted_data_buf[354] : n5194;   // modexp_top.v(481)
    assign n5203 = n2527 ? encrypted_data_buf[353] : n5195;   // modexp_top.v(481)
    assign n5204 = n2527 ? encrypted_data_buf[352] : n5196;   // modexp_top.v(481)
    assign n5205 = n2521 ? encrypted_data_buf[351] : n5197;   // modexp_top.v(481)
    assign n5206 = n2521 ? encrypted_data_buf[350] : n5198;   // modexp_top.v(481)
    assign n5207 = n2521 ? encrypted_data_buf[349] : n5199;   // modexp_top.v(481)
    assign n5208 = n2521 ? encrypted_data_buf[348] : n5200;   // modexp_top.v(481)
    assign n5209 = n2521 ? encrypted_data_buf[347] : n5201;   // modexp_top.v(481)
    assign n5210 = n2521 ? encrypted_data_buf[346] : n5202;   // modexp_top.v(481)
    assign n5211 = n2521 ? encrypted_data_buf[345] : n5203;   // modexp_top.v(481)
    assign n5212 = n2521 ? encrypted_data_buf[344] : n5204;   // modexp_top.v(481)
    assign n5213 = n2516 ? encrypted_data_buf[343] : n5205;   // modexp_top.v(481)
    assign n5214 = n2516 ? encrypted_data_buf[342] : n5206;   // modexp_top.v(481)
    assign n5215 = n2516 ? encrypted_data_buf[341] : n5207;   // modexp_top.v(481)
    assign n5216 = n2516 ? encrypted_data_buf[340] : n5208;   // modexp_top.v(481)
    assign n5217 = n2516 ? encrypted_data_buf[339] : n5209;   // modexp_top.v(481)
    assign n5218 = n2516 ? encrypted_data_buf[338] : n5210;   // modexp_top.v(481)
    assign n5219 = n2516 ? encrypted_data_buf[337] : n5211;   // modexp_top.v(481)
    assign n5220 = n2516 ? encrypted_data_buf[336] : n5212;   // modexp_top.v(481)
    assign n5221 = n2510 ? encrypted_data_buf[335] : n5213;   // modexp_top.v(481)
    assign n5222 = n2510 ? encrypted_data_buf[334] : n5214;   // modexp_top.v(481)
    assign n5223 = n2510 ? encrypted_data_buf[333] : n5215;   // modexp_top.v(481)
    assign n5224 = n2510 ? encrypted_data_buf[332] : n5216;   // modexp_top.v(481)
    assign n5225 = n2510 ? encrypted_data_buf[331] : n5217;   // modexp_top.v(481)
    assign n5226 = n2510 ? encrypted_data_buf[330] : n5218;   // modexp_top.v(481)
    assign n5227 = n2510 ? encrypted_data_buf[329] : n5219;   // modexp_top.v(481)
    assign n5228 = n2510 ? encrypted_data_buf[328] : n5220;   // modexp_top.v(481)
    assign n5229 = n2504 ? encrypted_data_buf[327] : n5221;   // modexp_top.v(481)
    assign n5230 = n2504 ? encrypted_data_buf[326] : n5222;   // modexp_top.v(481)
    assign n5231 = n2504 ? encrypted_data_buf[325] : n5223;   // modexp_top.v(481)
    assign n5232 = n2504 ? encrypted_data_buf[324] : n5224;   // modexp_top.v(481)
    assign n5233 = n2504 ? encrypted_data_buf[323] : n5225;   // modexp_top.v(481)
    assign n5234 = n2504 ? encrypted_data_buf[322] : n5226;   // modexp_top.v(481)
    assign n5235 = n2504 ? encrypted_data_buf[321] : n5227;   // modexp_top.v(481)
    assign n5236 = n2504 ? encrypted_data_buf[320] : n5228;   // modexp_top.v(481)
    assign n5237 = n2497 ? encrypted_data_buf[319] : n5229;   // modexp_top.v(481)
    assign n5238 = n2497 ? encrypted_data_buf[318] : n5230;   // modexp_top.v(481)
    assign n5239 = n2497 ? encrypted_data_buf[317] : n5231;   // modexp_top.v(481)
    assign n5240 = n2497 ? encrypted_data_buf[316] : n5232;   // modexp_top.v(481)
    assign n5241 = n2497 ? encrypted_data_buf[315] : n5233;   // modexp_top.v(481)
    assign n5242 = n2497 ? encrypted_data_buf[314] : n5234;   // modexp_top.v(481)
    assign n5243 = n2497 ? encrypted_data_buf[313] : n5235;   // modexp_top.v(481)
    assign n5244 = n2497 ? encrypted_data_buf[312] : n5236;   // modexp_top.v(481)
    assign n5245 = n2492 ? encrypted_data_buf[311] : n5237;   // modexp_top.v(481)
    assign n5246 = n2492 ? encrypted_data_buf[310] : n5238;   // modexp_top.v(481)
    assign n5247 = n2492 ? encrypted_data_buf[309] : n5239;   // modexp_top.v(481)
    assign n5248 = n2492 ? encrypted_data_buf[308] : n5240;   // modexp_top.v(481)
    assign n5249 = n2492 ? encrypted_data_buf[307] : n5241;   // modexp_top.v(481)
    assign n5250 = n2492 ? encrypted_data_buf[306] : n5242;   // modexp_top.v(481)
    assign n5251 = n2492 ? encrypted_data_buf[305] : n5243;   // modexp_top.v(481)
    assign n5252 = n2492 ? encrypted_data_buf[304] : n5244;   // modexp_top.v(481)
    assign n5253 = n2486 ? encrypted_data_buf[303] : n5245;   // modexp_top.v(481)
    assign n5254 = n2486 ? encrypted_data_buf[302] : n5246;   // modexp_top.v(481)
    assign n5255 = n2486 ? encrypted_data_buf[301] : n5247;   // modexp_top.v(481)
    assign n5256 = n2486 ? encrypted_data_buf[300] : n5248;   // modexp_top.v(481)
    assign n5257 = n2486 ? encrypted_data_buf[299] : n5249;   // modexp_top.v(481)
    assign n5258 = n2486 ? encrypted_data_buf[298] : n5250;   // modexp_top.v(481)
    assign n5259 = n2486 ? encrypted_data_buf[297] : n5251;   // modexp_top.v(481)
    assign n5260 = n2486 ? encrypted_data_buf[296] : n5252;   // modexp_top.v(481)
    assign n5261 = n2480 ? encrypted_data_buf[295] : n5253;   // modexp_top.v(481)
    assign n5262 = n2480 ? encrypted_data_buf[294] : n5254;   // modexp_top.v(481)
    assign n5263 = n2480 ? encrypted_data_buf[293] : n5255;   // modexp_top.v(481)
    assign n5264 = n2480 ? encrypted_data_buf[292] : n5256;   // modexp_top.v(481)
    assign n5265 = n2480 ? encrypted_data_buf[291] : n5257;   // modexp_top.v(481)
    assign n5266 = n2480 ? encrypted_data_buf[290] : n5258;   // modexp_top.v(481)
    assign n5267 = n2480 ? encrypted_data_buf[289] : n5259;   // modexp_top.v(481)
    assign n5268 = n2480 ? encrypted_data_buf[288] : n5260;   // modexp_top.v(481)
    assign n5269 = n2473 ? encrypted_data_buf[287] : n5261;   // modexp_top.v(481)
    assign n5270 = n2473 ? encrypted_data_buf[286] : n5262;   // modexp_top.v(481)
    assign n5271 = n2473 ? encrypted_data_buf[285] : n5263;   // modexp_top.v(481)
    assign n5272 = n2473 ? encrypted_data_buf[284] : n5264;   // modexp_top.v(481)
    assign n5273 = n2473 ? encrypted_data_buf[283] : n5265;   // modexp_top.v(481)
    assign n5274 = n2473 ? encrypted_data_buf[282] : n5266;   // modexp_top.v(481)
    assign n5275 = n2473 ? encrypted_data_buf[281] : n5267;   // modexp_top.v(481)
    assign n5276 = n2473 ? encrypted_data_buf[280] : n5268;   // modexp_top.v(481)
    assign n5277 = n2467 ? encrypted_data_buf[279] : n5269;   // modexp_top.v(481)
    assign n5278 = n2467 ? encrypted_data_buf[278] : n5270;   // modexp_top.v(481)
    assign n5279 = n2467 ? encrypted_data_buf[277] : n5271;   // modexp_top.v(481)
    assign n5280 = n2467 ? encrypted_data_buf[276] : n5272;   // modexp_top.v(481)
    assign n5281 = n2467 ? encrypted_data_buf[275] : n5273;   // modexp_top.v(481)
    assign n5282 = n2467 ? encrypted_data_buf[274] : n5274;   // modexp_top.v(481)
    assign n5283 = n2467 ? encrypted_data_buf[273] : n5275;   // modexp_top.v(481)
    assign n5284 = n2467 ? encrypted_data_buf[272] : n5276;   // modexp_top.v(481)
    assign n5285 = n2460 ? encrypted_data_buf[271] : n5277;   // modexp_top.v(481)
    assign n5286 = n2460 ? encrypted_data_buf[270] : n5278;   // modexp_top.v(481)
    assign n5287 = n2460 ? encrypted_data_buf[269] : n5279;   // modexp_top.v(481)
    assign n5288 = n2460 ? encrypted_data_buf[268] : n5280;   // modexp_top.v(481)
    assign n5289 = n2460 ? encrypted_data_buf[267] : n5281;   // modexp_top.v(481)
    assign n5290 = n2460 ? encrypted_data_buf[266] : n5282;   // modexp_top.v(481)
    assign n5291 = n2460 ? encrypted_data_buf[265] : n5283;   // modexp_top.v(481)
    assign n5292 = n2460 ? encrypted_data_buf[264] : n5284;   // modexp_top.v(481)
    assign n5293 = n2453 ? encrypted_data_buf[263] : n5285;   // modexp_top.v(481)
    assign n5294 = n2453 ? encrypted_data_buf[262] : n5286;   // modexp_top.v(481)
    assign n5295 = n2453 ? encrypted_data_buf[261] : n5287;   // modexp_top.v(481)
    assign n5296 = n2453 ? encrypted_data_buf[260] : n5288;   // modexp_top.v(481)
    assign n5297 = n2453 ? encrypted_data_buf[259] : n5289;   // modexp_top.v(481)
    assign n5298 = n2453 ? encrypted_data_buf[258] : n5290;   // modexp_top.v(481)
    assign n5299 = n2453 ? encrypted_data_buf[257] : n5291;   // modexp_top.v(481)
    assign n5300 = n2453 ? encrypted_data_buf[256] : n5292;   // modexp_top.v(481)
    assign n5301 = n2445 ? encrypted_data_buf[255] : n5293;   // modexp_top.v(481)
    assign n5302 = n2445 ? encrypted_data_buf[254] : n5294;   // modexp_top.v(481)
    assign n5303 = n2445 ? encrypted_data_buf[253] : n5295;   // modexp_top.v(481)
    assign n5304 = n2445 ? encrypted_data_buf[252] : n5296;   // modexp_top.v(481)
    assign n5305 = n2445 ? encrypted_data_buf[251] : n5297;   // modexp_top.v(481)
    assign n5306 = n2445 ? encrypted_data_buf[250] : n5298;   // modexp_top.v(481)
    assign n5307 = n2445 ? encrypted_data_buf[249] : n5299;   // modexp_top.v(481)
    assign n5308 = n2445 ? encrypted_data_buf[248] : n5300;   // modexp_top.v(481)
    assign n5309 = n2441 ? encrypted_data_buf[247] : n5301;   // modexp_top.v(481)
    assign n5310 = n2441 ? encrypted_data_buf[246] : n5302;   // modexp_top.v(481)
    assign n5311 = n2441 ? encrypted_data_buf[245] : n5303;   // modexp_top.v(481)
    assign n5312 = n2441 ? encrypted_data_buf[244] : n5304;   // modexp_top.v(481)
    assign n5313 = n2441 ? encrypted_data_buf[243] : n5305;   // modexp_top.v(481)
    assign n5314 = n2441 ? encrypted_data_buf[242] : n5306;   // modexp_top.v(481)
    assign n5315 = n2441 ? encrypted_data_buf[241] : n5307;   // modexp_top.v(481)
    assign n5316 = n2441 ? encrypted_data_buf[240] : n5308;   // modexp_top.v(481)
    assign n5317 = n2436 ? encrypted_data_buf[239] : n5309;   // modexp_top.v(481)
    assign n5318 = n2436 ? encrypted_data_buf[238] : n5310;   // modexp_top.v(481)
    assign n5319 = n2436 ? encrypted_data_buf[237] : n5311;   // modexp_top.v(481)
    assign n5320 = n2436 ? encrypted_data_buf[236] : n5312;   // modexp_top.v(481)
    assign n5321 = n2436 ? encrypted_data_buf[235] : n5313;   // modexp_top.v(481)
    assign n5322 = n2436 ? encrypted_data_buf[234] : n5314;   // modexp_top.v(481)
    assign n5323 = n2436 ? encrypted_data_buf[233] : n5315;   // modexp_top.v(481)
    assign n5324 = n2436 ? encrypted_data_buf[232] : n5316;   // modexp_top.v(481)
    assign n5325 = n2431 ? encrypted_data_buf[231] : n5317;   // modexp_top.v(481)
    assign n5326 = n2431 ? encrypted_data_buf[230] : n5318;   // modexp_top.v(481)
    assign n5327 = n2431 ? encrypted_data_buf[229] : n5319;   // modexp_top.v(481)
    assign n5328 = n2431 ? encrypted_data_buf[228] : n5320;   // modexp_top.v(481)
    assign n5329 = n2431 ? encrypted_data_buf[227] : n5321;   // modexp_top.v(481)
    assign n5330 = n2431 ? encrypted_data_buf[226] : n5322;   // modexp_top.v(481)
    assign n5331 = n2431 ? encrypted_data_buf[225] : n5323;   // modexp_top.v(481)
    assign n5332 = n2431 ? encrypted_data_buf[224] : n5324;   // modexp_top.v(481)
    assign n5333 = n2425 ? encrypted_data_buf[223] : n5325;   // modexp_top.v(481)
    assign n5334 = n2425 ? encrypted_data_buf[222] : n5326;   // modexp_top.v(481)
    assign n5335 = n2425 ? encrypted_data_buf[221] : n5327;   // modexp_top.v(481)
    assign n5336 = n2425 ? encrypted_data_buf[220] : n5328;   // modexp_top.v(481)
    assign n5337 = n2425 ? encrypted_data_buf[219] : n5329;   // modexp_top.v(481)
    assign n5338 = n2425 ? encrypted_data_buf[218] : n5330;   // modexp_top.v(481)
    assign n5339 = n2425 ? encrypted_data_buf[217] : n5331;   // modexp_top.v(481)
    assign n5340 = n2425 ? encrypted_data_buf[216] : n5332;   // modexp_top.v(481)
    assign n5341 = n2420 ? encrypted_data_buf[215] : n5333;   // modexp_top.v(481)
    assign n5342 = n2420 ? encrypted_data_buf[214] : n5334;   // modexp_top.v(481)
    assign n5343 = n2420 ? encrypted_data_buf[213] : n5335;   // modexp_top.v(481)
    assign n5344 = n2420 ? encrypted_data_buf[212] : n5336;   // modexp_top.v(481)
    assign n5345 = n2420 ? encrypted_data_buf[211] : n5337;   // modexp_top.v(481)
    assign n5346 = n2420 ? encrypted_data_buf[210] : n5338;   // modexp_top.v(481)
    assign n5347 = n2420 ? encrypted_data_buf[209] : n5339;   // modexp_top.v(481)
    assign n5348 = n2420 ? encrypted_data_buf[208] : n5340;   // modexp_top.v(481)
    assign n5349 = n2414 ? encrypted_data_buf[207] : n5341;   // modexp_top.v(481)
    assign n5350 = n2414 ? encrypted_data_buf[206] : n5342;   // modexp_top.v(481)
    assign n5351 = n2414 ? encrypted_data_buf[205] : n5343;   // modexp_top.v(481)
    assign n5352 = n2414 ? encrypted_data_buf[204] : n5344;   // modexp_top.v(481)
    assign n5353 = n2414 ? encrypted_data_buf[203] : n5345;   // modexp_top.v(481)
    assign n5354 = n2414 ? encrypted_data_buf[202] : n5346;   // modexp_top.v(481)
    assign n5355 = n2414 ? encrypted_data_buf[201] : n5347;   // modexp_top.v(481)
    assign n5356 = n2414 ? encrypted_data_buf[200] : n5348;   // modexp_top.v(481)
    assign n5357 = n2408 ? encrypted_data_buf[199] : n5349;   // modexp_top.v(481)
    assign n5358 = n2408 ? encrypted_data_buf[198] : n5350;   // modexp_top.v(481)
    assign n5359 = n2408 ? encrypted_data_buf[197] : n5351;   // modexp_top.v(481)
    assign n5360 = n2408 ? encrypted_data_buf[196] : n5352;   // modexp_top.v(481)
    assign n5361 = n2408 ? encrypted_data_buf[195] : n5353;   // modexp_top.v(481)
    assign n5362 = n2408 ? encrypted_data_buf[194] : n5354;   // modexp_top.v(481)
    assign n5363 = n2408 ? encrypted_data_buf[193] : n5355;   // modexp_top.v(481)
    assign n5364 = n2408 ? encrypted_data_buf[192] : n5356;   // modexp_top.v(481)
    assign n5365 = n2401 ? encrypted_data_buf[191] : n5357;   // modexp_top.v(481)
    assign n5366 = n2401 ? encrypted_data_buf[190] : n5358;   // modexp_top.v(481)
    assign n5367 = n2401 ? encrypted_data_buf[189] : n5359;   // modexp_top.v(481)
    assign n5368 = n2401 ? encrypted_data_buf[188] : n5360;   // modexp_top.v(481)
    assign n5369 = n2401 ? encrypted_data_buf[187] : n5361;   // modexp_top.v(481)
    assign n5370 = n2401 ? encrypted_data_buf[186] : n5362;   // modexp_top.v(481)
    assign n5371 = n2401 ? encrypted_data_buf[185] : n5363;   // modexp_top.v(481)
    assign n5372 = n2401 ? encrypted_data_buf[184] : n5364;   // modexp_top.v(481)
    assign n5373 = n2396 ? encrypted_data_buf[183] : n5365;   // modexp_top.v(481)
    assign n5374 = n2396 ? encrypted_data_buf[182] : n5366;   // modexp_top.v(481)
    assign n5375 = n2396 ? encrypted_data_buf[181] : n5367;   // modexp_top.v(481)
    assign n5376 = n2396 ? encrypted_data_buf[180] : n5368;   // modexp_top.v(481)
    assign n5377 = n2396 ? encrypted_data_buf[179] : n5369;   // modexp_top.v(481)
    assign n5378 = n2396 ? encrypted_data_buf[178] : n5370;   // modexp_top.v(481)
    assign n5379 = n2396 ? encrypted_data_buf[177] : n5371;   // modexp_top.v(481)
    assign n5380 = n2396 ? encrypted_data_buf[176] : n5372;   // modexp_top.v(481)
    assign n5381 = n2390 ? encrypted_data_buf[175] : n5373;   // modexp_top.v(481)
    assign n5382 = n2390 ? encrypted_data_buf[174] : n5374;   // modexp_top.v(481)
    assign n5383 = n2390 ? encrypted_data_buf[173] : n5375;   // modexp_top.v(481)
    assign n5384 = n2390 ? encrypted_data_buf[172] : n5376;   // modexp_top.v(481)
    assign n5385 = n2390 ? encrypted_data_buf[171] : n5377;   // modexp_top.v(481)
    assign n5386 = n2390 ? encrypted_data_buf[170] : n5378;   // modexp_top.v(481)
    assign n5387 = n2390 ? encrypted_data_buf[169] : n5379;   // modexp_top.v(481)
    assign n5388 = n2390 ? encrypted_data_buf[168] : n5380;   // modexp_top.v(481)
    assign n5389 = n2384 ? encrypted_data_buf[167] : n5381;   // modexp_top.v(481)
    assign n5390 = n2384 ? encrypted_data_buf[166] : n5382;   // modexp_top.v(481)
    assign n5391 = n2384 ? encrypted_data_buf[165] : n5383;   // modexp_top.v(481)
    assign n5392 = n2384 ? encrypted_data_buf[164] : n5384;   // modexp_top.v(481)
    assign n5393 = n2384 ? encrypted_data_buf[163] : n5385;   // modexp_top.v(481)
    assign n5394 = n2384 ? encrypted_data_buf[162] : n5386;   // modexp_top.v(481)
    assign n5395 = n2384 ? encrypted_data_buf[161] : n5387;   // modexp_top.v(481)
    assign n5396 = n2384 ? encrypted_data_buf[160] : n5388;   // modexp_top.v(481)
    assign n5397 = n2377 ? encrypted_data_buf[159] : n5389;   // modexp_top.v(481)
    assign n5398 = n2377 ? encrypted_data_buf[158] : n5390;   // modexp_top.v(481)
    assign n5399 = n2377 ? encrypted_data_buf[157] : n5391;   // modexp_top.v(481)
    assign n5400 = n2377 ? encrypted_data_buf[156] : n5392;   // modexp_top.v(481)
    assign n5401 = n2377 ? encrypted_data_buf[155] : n5393;   // modexp_top.v(481)
    assign n5402 = n2377 ? encrypted_data_buf[154] : n5394;   // modexp_top.v(481)
    assign n5403 = n2377 ? encrypted_data_buf[153] : n5395;   // modexp_top.v(481)
    assign n5404 = n2377 ? encrypted_data_buf[152] : n5396;   // modexp_top.v(481)
    assign n5405 = n2371 ? encrypted_data_buf[151] : n5397;   // modexp_top.v(481)
    assign n5406 = n2371 ? encrypted_data_buf[150] : n5398;   // modexp_top.v(481)
    assign n5407 = n2371 ? encrypted_data_buf[149] : n5399;   // modexp_top.v(481)
    assign n5408 = n2371 ? encrypted_data_buf[148] : n5400;   // modexp_top.v(481)
    assign n5409 = n2371 ? encrypted_data_buf[147] : n5401;   // modexp_top.v(481)
    assign n5410 = n2371 ? encrypted_data_buf[146] : n5402;   // modexp_top.v(481)
    assign n5411 = n2371 ? encrypted_data_buf[145] : n5403;   // modexp_top.v(481)
    assign n5412 = n2371 ? encrypted_data_buf[144] : n5404;   // modexp_top.v(481)
    assign n5413 = n2364 ? encrypted_data_buf[143] : n5405;   // modexp_top.v(481)
    assign n5414 = n2364 ? encrypted_data_buf[142] : n5406;   // modexp_top.v(481)
    assign n5415 = n2364 ? encrypted_data_buf[141] : n5407;   // modexp_top.v(481)
    assign n5416 = n2364 ? encrypted_data_buf[140] : n5408;   // modexp_top.v(481)
    assign n5417 = n2364 ? encrypted_data_buf[139] : n5409;   // modexp_top.v(481)
    assign n5418 = n2364 ? encrypted_data_buf[138] : n5410;   // modexp_top.v(481)
    assign n5419 = n2364 ? encrypted_data_buf[137] : n5411;   // modexp_top.v(481)
    assign n5420 = n2364 ? encrypted_data_buf[136] : n5412;   // modexp_top.v(481)
    assign n5421 = n2357 ? encrypted_data_buf[135] : n5413;   // modexp_top.v(481)
    assign n5422 = n2357 ? encrypted_data_buf[134] : n5414;   // modexp_top.v(481)
    assign n5423 = n2357 ? encrypted_data_buf[133] : n5415;   // modexp_top.v(481)
    assign n5424 = n2357 ? encrypted_data_buf[132] : n5416;   // modexp_top.v(481)
    assign n5425 = n2357 ? encrypted_data_buf[131] : n5417;   // modexp_top.v(481)
    assign n5426 = n2357 ? encrypted_data_buf[130] : n5418;   // modexp_top.v(481)
    assign n5427 = n2357 ? encrypted_data_buf[129] : n5419;   // modexp_top.v(481)
    assign n5428 = n2357 ? encrypted_data_buf[128] : n5420;   // modexp_top.v(481)
    assign n5429 = n2349 ? encrypted_data_buf[127] : n5421;   // modexp_top.v(481)
    assign n5430 = n2349 ? encrypted_data_buf[126] : n5422;   // modexp_top.v(481)
    assign n5431 = n2349 ? encrypted_data_buf[125] : n5423;   // modexp_top.v(481)
    assign n5432 = n2349 ? encrypted_data_buf[124] : n5424;   // modexp_top.v(481)
    assign n5433 = n2349 ? encrypted_data_buf[123] : n5425;   // modexp_top.v(481)
    assign n5434 = n2349 ? encrypted_data_buf[122] : n5426;   // modexp_top.v(481)
    assign n5435 = n2349 ? encrypted_data_buf[121] : n5427;   // modexp_top.v(481)
    assign n5436 = n2349 ? encrypted_data_buf[120] : n5428;   // modexp_top.v(481)
    assign n5437 = n2344 ? encrypted_data_buf[119] : n5429;   // modexp_top.v(481)
    assign n5438 = n2344 ? encrypted_data_buf[118] : n5430;   // modexp_top.v(481)
    assign n5439 = n2344 ? encrypted_data_buf[117] : n5431;   // modexp_top.v(481)
    assign n5440 = n2344 ? encrypted_data_buf[116] : n5432;   // modexp_top.v(481)
    assign n5441 = n2344 ? encrypted_data_buf[115] : n5433;   // modexp_top.v(481)
    assign n5442 = n2344 ? encrypted_data_buf[114] : n5434;   // modexp_top.v(481)
    assign n5443 = n2344 ? encrypted_data_buf[113] : n5435;   // modexp_top.v(481)
    assign n5444 = n2344 ? encrypted_data_buf[112] : n5436;   // modexp_top.v(481)
    assign n5445 = n2338 ? encrypted_data_buf[111] : n5437;   // modexp_top.v(481)
    assign n5446 = n2338 ? encrypted_data_buf[110] : n5438;   // modexp_top.v(481)
    assign n5447 = n2338 ? encrypted_data_buf[109] : n5439;   // modexp_top.v(481)
    assign n5448 = n2338 ? encrypted_data_buf[108] : n5440;   // modexp_top.v(481)
    assign n5449 = n2338 ? encrypted_data_buf[107] : n5441;   // modexp_top.v(481)
    assign n5450 = n2338 ? encrypted_data_buf[106] : n5442;   // modexp_top.v(481)
    assign n5451 = n2338 ? encrypted_data_buf[105] : n5443;   // modexp_top.v(481)
    assign n5452 = n2338 ? encrypted_data_buf[104] : n5444;   // modexp_top.v(481)
    assign n5453 = n2332 ? encrypted_data_buf[103] : n5445;   // modexp_top.v(481)
    assign n5454 = n2332 ? encrypted_data_buf[102] : n5446;   // modexp_top.v(481)
    assign n5455 = n2332 ? encrypted_data_buf[101] : n5447;   // modexp_top.v(481)
    assign n5456 = n2332 ? encrypted_data_buf[100] : n5448;   // modexp_top.v(481)
    assign n5457 = n2332 ? encrypted_data_buf[99] : n5449;   // modexp_top.v(481)
    assign n5458 = n2332 ? encrypted_data_buf[98] : n5450;   // modexp_top.v(481)
    assign n5459 = n2332 ? encrypted_data_buf[97] : n5451;   // modexp_top.v(481)
    assign n5460 = n2332 ? encrypted_data_buf[96] : n5452;   // modexp_top.v(481)
    assign n5461 = n2325 ? encrypted_data_buf[95] : n5453;   // modexp_top.v(481)
    assign n5462 = n2325 ? encrypted_data_buf[94] : n5454;   // modexp_top.v(481)
    assign n5463 = n2325 ? encrypted_data_buf[93] : n5455;   // modexp_top.v(481)
    assign n5464 = n2325 ? encrypted_data_buf[92] : n5456;   // modexp_top.v(481)
    assign n5465 = n2325 ? encrypted_data_buf[91] : n5457;   // modexp_top.v(481)
    assign n5466 = n2325 ? encrypted_data_buf[90] : n5458;   // modexp_top.v(481)
    assign n5467 = n2325 ? encrypted_data_buf[89] : n5459;   // modexp_top.v(481)
    assign n5468 = n2325 ? encrypted_data_buf[88] : n5460;   // modexp_top.v(481)
    assign n5469 = n2319 ? encrypted_data_buf[87] : n5461;   // modexp_top.v(481)
    assign n5470 = n2319 ? encrypted_data_buf[86] : n5462;   // modexp_top.v(481)
    assign n5471 = n2319 ? encrypted_data_buf[85] : n5463;   // modexp_top.v(481)
    assign n5472 = n2319 ? encrypted_data_buf[84] : n5464;   // modexp_top.v(481)
    assign n5473 = n2319 ? encrypted_data_buf[83] : n5465;   // modexp_top.v(481)
    assign n5474 = n2319 ? encrypted_data_buf[82] : n5466;   // modexp_top.v(481)
    assign n5475 = n2319 ? encrypted_data_buf[81] : n5467;   // modexp_top.v(481)
    assign n5476 = n2319 ? encrypted_data_buf[80] : n5468;   // modexp_top.v(481)
    assign n5477 = n2312 ? encrypted_data_buf[79] : n5469;   // modexp_top.v(481)
    assign n5478 = n2312 ? encrypted_data_buf[78] : n5470;   // modexp_top.v(481)
    assign n5479 = n2312 ? encrypted_data_buf[77] : n5471;   // modexp_top.v(481)
    assign n5480 = n2312 ? encrypted_data_buf[76] : n5472;   // modexp_top.v(481)
    assign n5481 = n2312 ? encrypted_data_buf[75] : n5473;   // modexp_top.v(481)
    assign n5482 = n2312 ? encrypted_data_buf[74] : n5474;   // modexp_top.v(481)
    assign n5483 = n2312 ? encrypted_data_buf[73] : n5475;   // modexp_top.v(481)
    assign n5484 = n2312 ? encrypted_data_buf[72] : n5476;   // modexp_top.v(481)
    assign n5485 = n2305 ? encrypted_data_buf[71] : n5477;   // modexp_top.v(481)
    assign n5486 = n2305 ? encrypted_data_buf[70] : n5478;   // modexp_top.v(481)
    assign n5487 = n2305 ? encrypted_data_buf[69] : n5479;   // modexp_top.v(481)
    assign n5488 = n2305 ? encrypted_data_buf[68] : n5480;   // modexp_top.v(481)
    assign n5489 = n2305 ? encrypted_data_buf[67] : n5481;   // modexp_top.v(481)
    assign n5490 = n2305 ? encrypted_data_buf[66] : n5482;   // modexp_top.v(481)
    assign n5491 = n2305 ? encrypted_data_buf[65] : n5483;   // modexp_top.v(481)
    assign n5492 = n2305 ? encrypted_data_buf[64] : n5484;   // modexp_top.v(481)
    assign n5493 = n2297 ? encrypted_data_buf[63] : n5485;   // modexp_top.v(481)
    assign n5494 = n2297 ? encrypted_data_buf[62] : n5486;   // modexp_top.v(481)
    assign n5495 = n2297 ? encrypted_data_buf[61] : n5487;   // modexp_top.v(481)
    assign n5496 = n2297 ? encrypted_data_buf[60] : n5488;   // modexp_top.v(481)
    assign n5497 = n2297 ? encrypted_data_buf[59] : n5489;   // modexp_top.v(481)
    assign n5498 = n2297 ? encrypted_data_buf[58] : n5490;   // modexp_top.v(481)
    assign n5499 = n2297 ? encrypted_data_buf[57] : n5491;   // modexp_top.v(481)
    assign n5500 = n2297 ? encrypted_data_buf[56] : n5492;   // modexp_top.v(481)
    assign n5501 = n2291 ? encrypted_data_buf[55] : n5493;   // modexp_top.v(481)
    assign n5502 = n2291 ? encrypted_data_buf[54] : n5494;   // modexp_top.v(481)
    assign n5503 = n2291 ? encrypted_data_buf[53] : n5495;   // modexp_top.v(481)
    assign n5504 = n2291 ? encrypted_data_buf[52] : n5496;   // modexp_top.v(481)
    assign n5505 = n2291 ? encrypted_data_buf[51] : n5497;   // modexp_top.v(481)
    assign n5506 = n2291 ? encrypted_data_buf[50] : n5498;   // modexp_top.v(481)
    assign n5507 = n2291 ? encrypted_data_buf[49] : n5499;   // modexp_top.v(481)
    assign n5508 = n2291 ? encrypted_data_buf[48] : n5500;   // modexp_top.v(481)
    assign n5509 = n2284 ? encrypted_data_buf[47] : n5501;   // modexp_top.v(481)
    assign n5510 = n2284 ? encrypted_data_buf[46] : n5502;   // modexp_top.v(481)
    assign n5511 = n2284 ? encrypted_data_buf[45] : n5503;   // modexp_top.v(481)
    assign n5512 = n2284 ? encrypted_data_buf[44] : n5504;   // modexp_top.v(481)
    assign n5513 = n2284 ? encrypted_data_buf[43] : n5505;   // modexp_top.v(481)
    assign n5514 = n2284 ? encrypted_data_buf[42] : n5506;   // modexp_top.v(481)
    assign n5515 = n2284 ? encrypted_data_buf[41] : n5507;   // modexp_top.v(481)
    assign n5516 = n2284 ? encrypted_data_buf[40] : n5508;   // modexp_top.v(481)
    assign n5517 = n2277 ? encrypted_data_buf[39] : n5509;   // modexp_top.v(481)
    assign n5518 = n2277 ? encrypted_data_buf[38] : n5510;   // modexp_top.v(481)
    assign n5519 = n2277 ? encrypted_data_buf[37] : n5511;   // modexp_top.v(481)
    assign n5520 = n2277 ? encrypted_data_buf[36] : n5512;   // modexp_top.v(481)
    assign n5521 = n2277 ? encrypted_data_buf[35] : n5513;   // modexp_top.v(481)
    assign n5522 = n2277 ? encrypted_data_buf[34] : n5514;   // modexp_top.v(481)
    assign n5523 = n2277 ? encrypted_data_buf[33] : n5515;   // modexp_top.v(481)
    assign n5524 = n2277 ? encrypted_data_buf[32] : n5516;   // modexp_top.v(481)
    assign n5525 = n2269 ? encrypted_data_buf[31] : n5517;   // modexp_top.v(481)
    assign n5526 = n2269 ? encrypted_data_buf[30] : n5518;   // modexp_top.v(481)
    assign n5527 = n2269 ? encrypted_data_buf[29] : n5519;   // modexp_top.v(481)
    assign n5528 = n2269 ? encrypted_data_buf[28] : n5520;   // modexp_top.v(481)
    assign n5529 = n2269 ? encrypted_data_buf[27] : n5521;   // modexp_top.v(481)
    assign n5530 = n2269 ? encrypted_data_buf[26] : n5522;   // modexp_top.v(481)
    assign n5531 = n2269 ? encrypted_data_buf[25] : n5523;   // modexp_top.v(481)
    assign n5532 = n2269 ? encrypted_data_buf[24] : n5524;   // modexp_top.v(481)
    assign n5533 = n2262 ? encrypted_data_buf[23] : n5525;   // modexp_top.v(481)
    assign n5534 = n2262 ? encrypted_data_buf[22] : n5526;   // modexp_top.v(481)
    assign n5535 = n2262 ? encrypted_data_buf[21] : n5527;   // modexp_top.v(481)
    assign n5536 = n2262 ? encrypted_data_buf[20] : n5528;   // modexp_top.v(481)
    assign n5537 = n2262 ? encrypted_data_buf[19] : n5529;   // modexp_top.v(481)
    assign n5538 = n2262 ? encrypted_data_buf[18] : n5530;   // modexp_top.v(481)
    assign n5539 = n2262 ? encrypted_data_buf[17] : n5531;   // modexp_top.v(481)
    assign n5540 = n2262 ? encrypted_data_buf[16] : n5532;   // modexp_top.v(481)
    assign n5541 = n2254 ? encrypted_data_buf[15] : n5533;   // modexp_top.v(481)
    assign n5542 = n2254 ? encrypted_data_buf[14] : n5534;   // modexp_top.v(481)
    assign n5543 = n2254 ? encrypted_data_buf[13] : n5535;   // modexp_top.v(481)
    assign n5544 = n2254 ? encrypted_data_buf[12] : n5536;   // modexp_top.v(481)
    assign n5545 = n2254 ? encrypted_data_buf[11] : n5537;   // modexp_top.v(481)
    assign n5546 = n2254 ? encrypted_data_buf[10] : n5538;   // modexp_top.v(481)
    assign n5547 = n2254 ? encrypted_data_buf[9] : n5539;   // modexp_top.v(481)
    assign n5548 = n2254 ? encrypted_data_buf[8] : n5540;   // modexp_top.v(481)
    assign xram_data_out[7] = n2246 ? encrypted_data_buf[7] : n5541;   // modexp_top.v(481)
    assign xram_data_out[6] = n2246 ? encrypted_data_buf[6] : n5542;   // modexp_top.v(481)
    assign xram_data_out[5] = n2246 ? encrypted_data_buf[5] : n5543;   // modexp_top.v(481)
    assign xram_data_out[4] = n2246 ? encrypted_data_buf[4] : n5544;   // modexp_top.v(481)
    assign xram_data_out[3] = n2246 ? encrypted_data_buf[3] : n5545;   // modexp_top.v(481)
    assign xram_data_out[2] = n2246 ? encrypted_data_buf[2] : n5546;   // modexp_top.v(481)
    assign xram_data_out[1] = n2246 ? encrypted_data_buf[1] : n5547;   // modexp_top.v(481)
    assign xram_data_out[0] = n2246 ? encrypted_data_buf[0] : n5548;   // modexp_top.v(481)
    VERIFIC_DFFRS i5535 (.d(exp_reg_state_next[0]), .clk(clk), .s(1'b0), 
            .r(rst), .q(exp_state[0]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5536 (.d(byte_counter_next[7]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[7]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5537 (.d(byte_counter_next[6]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[6]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5538 (.d(byte_counter_next[5]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[5]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5539 (.d(byte_counter_next[4]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[4]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5540 (.d(byte_counter_next[3]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[3]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5541 (.d(byte_counter_next[2]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[2]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5542 (.d(byte_counter_next[1]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[1]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5543 (.d(byte_counter_next[0]), .clk(clk), .s(1'b0), 
            .r(rst), .q(byte_counter[0]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5544 (.d(n7616), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2047]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5545 (.d(n7617), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2046]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5546 (.d(n7618), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2045]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5547 (.d(n7619), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2044]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5548 (.d(n7620), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2043]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5549 (.d(n7621), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2042]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5550 (.d(n7622), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2041]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5551 (.d(n7623), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2040]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5552 (.d(n7624), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2039]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5553 (.d(n7625), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2038]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5554 (.d(n7626), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2037]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5555 (.d(n7627), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2036]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5556 (.d(n7628), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2035]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5557 (.d(n7629), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2034]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5558 (.d(n7630), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2033]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5559 (.d(n7631), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2032]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5560 (.d(n7632), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2031]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5561 (.d(n7633), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2030]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5562 (.d(n7634), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2029]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5563 (.d(n7635), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2028]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5564 (.d(n7636), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2027]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5565 (.d(n7637), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2026]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5566 (.d(n7638), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2025]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5567 (.d(n7639), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2024]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5568 (.d(n7640), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2023]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5569 (.d(n7641), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2022]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5570 (.d(n7642), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2021]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5571 (.d(n7643), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2020]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5572 (.d(n7644), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2019]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5573 (.d(n7645), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2018]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5574 (.d(n7646), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2017]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5575 (.d(n7647), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2016]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5576 (.d(n7648), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2015]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5577 (.d(n7649), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2014]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5578 (.d(n7650), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2013]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5579 (.d(n7651), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2012]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5580 (.d(n7652), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2011]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5581 (.d(n7653), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2010]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5582 (.d(n7654), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2009]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5583 (.d(n7655), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2008]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5584 (.d(n7656), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2007]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5585 (.d(n7657), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2006]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5586 (.d(n7658), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2005]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5587 (.d(n7659), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2004]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5588 (.d(n7660), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2003]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5589 (.d(n7661), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2002]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5590 (.d(n7662), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2001]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5591 (.d(n7663), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2000]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5592 (.d(n7664), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1999]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5593 (.d(n7665), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1998]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5594 (.d(n7666), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1997]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5595 (.d(n7667), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1996]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5596 (.d(n7668), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1995]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5597 (.d(n7669), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1994]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5598 (.d(n7670), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1993]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5599 (.d(n7671), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1992]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5600 (.d(n7672), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1991]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5601 (.d(n7673), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1990]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5602 (.d(n7674), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1989]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5603 (.d(n7675), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1988]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5604 (.d(n7676), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1987]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5605 (.d(n7677), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1986]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5606 (.d(n7678), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1985]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5607 (.d(n7679), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1984]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5608 (.d(n7680), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1983]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5609 (.d(n7681), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1982]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5610 (.d(n7682), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1981]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5611 (.d(n7683), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1980]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5612 (.d(n7684), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1979]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5613 (.d(n7685), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1978]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5614 (.d(n7686), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1977]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5615 (.d(n7687), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1976]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5616 (.d(n7688), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1975]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5617 (.d(n7689), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1974]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5618 (.d(n7690), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1973]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5619 (.d(n7691), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1972]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5620 (.d(n7692), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1971]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5621 (.d(n7693), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1970]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5622 (.d(n7694), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1969]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5623 (.d(n7695), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1968]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5624 (.d(n7696), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1967]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5625 (.d(n7697), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1966]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5626 (.d(n7698), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1965]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5627 (.d(n7699), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1964]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5628 (.d(n7700), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1963]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5629 (.d(n7701), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1962]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5630 (.d(n7702), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1961]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5631 (.d(n7703), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1960]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5632 (.d(n7704), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1959]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5633 (.d(n7705), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1958]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5634 (.d(n7706), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1957]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5635 (.d(n7707), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1956]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5636 (.d(n7708), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1955]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5637 (.d(n7709), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1954]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5638 (.d(n7710), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1953]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5639 (.d(n7711), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1952]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5640 (.d(n7712), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1951]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5641 (.d(n7713), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1950]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5642 (.d(n7714), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1949]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5643 (.d(n7715), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1948]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5644 (.d(n7716), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1947]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5645 (.d(n7717), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1946]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5646 (.d(n7718), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1945]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5647 (.d(n7719), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1944]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5648 (.d(n7720), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1943]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5649 (.d(n7721), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1942]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5650 (.d(n7722), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1941]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5651 (.d(n7723), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1940]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5652 (.d(n7724), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1939]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5653 (.d(n7725), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1938]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5654 (.d(n7726), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1937]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5655 (.d(n7727), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1936]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5656 (.d(n7728), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1935]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5657 (.d(n7729), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1934]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5658 (.d(n7730), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1933]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5659 (.d(n7731), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1932]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5660 (.d(n7732), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1931]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5661 (.d(n7733), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1930]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5662 (.d(n7734), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1929]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5663 (.d(n7735), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1928]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5664 (.d(n7736), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1927]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5665 (.d(n7737), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1926]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5666 (.d(n7738), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1925]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5667 (.d(n7739), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1924]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5668 (.d(n7740), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1923]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5669 (.d(n7741), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1922]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5670 (.d(n7742), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1921]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5671 (.d(n7743), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1920]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5672 (.d(n7744), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1919]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5673 (.d(n7745), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1918]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5674 (.d(n7746), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1917]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5675 (.d(n7747), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1916]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5676 (.d(n7748), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1915]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5677 (.d(n7749), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1914]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5678 (.d(n7750), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1913]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5679 (.d(n7751), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1912]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5680 (.d(n7752), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1911]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5681 (.d(n7753), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1910]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5682 (.d(n7754), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1909]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5683 (.d(n7755), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1908]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5684 (.d(n7756), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1907]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5685 (.d(n7757), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1906]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5686 (.d(n7758), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1905]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5687 (.d(n7759), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1904]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5688 (.d(n7760), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1903]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5689 (.d(n7761), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1902]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5690 (.d(n7762), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1901]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5691 (.d(n7763), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1900]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5692 (.d(n7764), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1899]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5693 (.d(n7765), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1898]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5694 (.d(n7766), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1897]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5695 (.d(n7767), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1896]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5696 (.d(n7768), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1895]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5697 (.d(n7769), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1894]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5698 (.d(n7770), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1893]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5699 (.d(n7771), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1892]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5700 (.d(n7772), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1891]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5701 (.d(n7773), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1890]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5702 (.d(n7774), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1889]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5703 (.d(n7775), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1888]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5704 (.d(n7776), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1887]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5705 (.d(n7777), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1886]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5706 (.d(n7778), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1885]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5707 (.d(n7779), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1884]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5708 (.d(n7780), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1883]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5709 (.d(n7781), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1882]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5710 (.d(n7782), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1881]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5711 (.d(n7783), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1880]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5712 (.d(n7784), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1879]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5713 (.d(n7785), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1878]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5714 (.d(n7786), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1877]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5715 (.d(n7787), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1876]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5716 (.d(n7788), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1875]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5717 (.d(n7789), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1874]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5718 (.d(n7790), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1873]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5719 (.d(n7791), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1872]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5720 (.d(n7792), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1871]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5721 (.d(n7793), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1870]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5722 (.d(n7794), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1869]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5723 (.d(n7795), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1868]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5724 (.d(n7796), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1867]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5725 (.d(n7797), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1866]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5726 (.d(n7798), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1865]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5727 (.d(n7799), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1864]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5728 (.d(n7800), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1863]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5729 (.d(n7801), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1862]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5730 (.d(n7802), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1861]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5731 (.d(n7803), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1860]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5732 (.d(n7804), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1859]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5733 (.d(n7805), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1858]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5734 (.d(n7806), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1857]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5735 (.d(n7807), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1856]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5736 (.d(n7808), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1855]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5737 (.d(n7809), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1854]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5738 (.d(n7810), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1853]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5739 (.d(n7811), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1852]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5740 (.d(n7812), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1851]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5741 (.d(n7813), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1850]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5742 (.d(n7814), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1849]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5743 (.d(n7815), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1848]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5744 (.d(n7816), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1847]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5745 (.d(n7817), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1846]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5746 (.d(n7818), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1845]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5747 (.d(n7819), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1844]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5748 (.d(n7820), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1843]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5749 (.d(n7821), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1842]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5750 (.d(n7822), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1841]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5751 (.d(n7823), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1840]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5752 (.d(n7824), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1839]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5753 (.d(n7825), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1838]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5754 (.d(n7826), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1837]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5755 (.d(n7827), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1836]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5756 (.d(n7828), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1835]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5757 (.d(n7829), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1834]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5758 (.d(n7830), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1833]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5759 (.d(n7831), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1832]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5760 (.d(n7832), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1831]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5761 (.d(n7833), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1830]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5762 (.d(n7834), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1829]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5763 (.d(n7835), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1828]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5764 (.d(n7836), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1827]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5765 (.d(n7837), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1826]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5766 (.d(n7838), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1825]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5767 (.d(n7839), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1824]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5768 (.d(n7840), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1823]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5769 (.d(n7841), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1822]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5770 (.d(n7842), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1821]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5771 (.d(n7843), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1820]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5772 (.d(n7844), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1819]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5773 (.d(n7845), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1818]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5774 (.d(n7846), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1817]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5775 (.d(n7847), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1816]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5776 (.d(n7848), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1815]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5777 (.d(n7849), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1814]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5778 (.d(n7850), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1813]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5779 (.d(n7851), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1812]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5780 (.d(n7852), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1811]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5781 (.d(n7853), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1810]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5782 (.d(n7854), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1809]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5783 (.d(n7855), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1808]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5784 (.d(n7856), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1807]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5785 (.d(n7857), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1806]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5786 (.d(n7858), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1805]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5787 (.d(n7859), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1804]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5788 (.d(n7860), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1803]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5789 (.d(n7861), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1802]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5790 (.d(n7862), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1801]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5791 (.d(n7863), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1800]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5792 (.d(n7864), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1799]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5793 (.d(n7865), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1798]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5794 (.d(n7866), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1797]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5795 (.d(n7867), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1796]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5796 (.d(n7868), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1795]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5797 (.d(n7869), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1794]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5798 (.d(n7870), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1793]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5799 (.d(n7871), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1792]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5800 (.d(n7872), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1791]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5801 (.d(n7873), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1790]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5802 (.d(n7874), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1789]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5803 (.d(n7875), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1788]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5804 (.d(n7876), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1787]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5805 (.d(n7877), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1786]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5806 (.d(n7878), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1785]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5807 (.d(n7879), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1784]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5808 (.d(n7880), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1783]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5809 (.d(n7881), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1782]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5810 (.d(n7882), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1781]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5811 (.d(n7883), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1780]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5812 (.d(n7884), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1779]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5813 (.d(n7885), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1778]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5814 (.d(n7886), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1777]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5815 (.d(n7887), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1776]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5816 (.d(n7888), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1775]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5817 (.d(n7889), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1774]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5818 (.d(n7890), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1773]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5819 (.d(n7891), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1772]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5820 (.d(n7892), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1771]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5821 (.d(n7893), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1770]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5822 (.d(n7894), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1769]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5823 (.d(n7895), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1768]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5824 (.d(n7896), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1767]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5825 (.d(n7897), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1766]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5826 (.d(n7898), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1765]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5827 (.d(n7899), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1764]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5828 (.d(n7900), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1763]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5829 (.d(n7901), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1762]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5830 (.d(n7902), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1761]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5831 (.d(n7903), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1760]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5832 (.d(n7904), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1759]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5833 (.d(n7905), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1758]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5834 (.d(n7906), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1757]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5835 (.d(n7907), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1756]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5836 (.d(n7908), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1755]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5837 (.d(n7909), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1754]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5838 (.d(n7910), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1753]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5839 (.d(n7911), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1752]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5840 (.d(n7912), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1751]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5841 (.d(n7913), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1750]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5842 (.d(n7914), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1749]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5843 (.d(n7915), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1748]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5844 (.d(n7916), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1747]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5845 (.d(n7917), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1746]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5846 (.d(n7918), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1745]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5847 (.d(n7919), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1744]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5848 (.d(n7920), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1743]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5849 (.d(n7921), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1742]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5850 (.d(n7922), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1741]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5851 (.d(n7923), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1740]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5852 (.d(n7924), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1739]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5853 (.d(n7925), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1738]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5854 (.d(n7926), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1737]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5855 (.d(n7927), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1736]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5856 (.d(n7928), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1735]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5857 (.d(n7929), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1734]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5858 (.d(n7930), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1733]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5859 (.d(n7931), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1732]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5860 (.d(n7932), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1731]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5861 (.d(n7933), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1730]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5862 (.d(n7934), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1729]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5863 (.d(n7935), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1728]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5864 (.d(n7936), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1727]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5865 (.d(n7937), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1726]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5866 (.d(n7938), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1725]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5867 (.d(n7939), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1724]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5868 (.d(n7940), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1723]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5869 (.d(n7941), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1722]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5870 (.d(n7942), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1721]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5871 (.d(n7943), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1720]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5872 (.d(n7944), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1719]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5873 (.d(n7945), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1718]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5874 (.d(n7946), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1717]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5875 (.d(n7947), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1716]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5876 (.d(n7948), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1715]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5877 (.d(n7949), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1714]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5878 (.d(n7950), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1713]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5879 (.d(n7951), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1712]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5880 (.d(n7952), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1711]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5881 (.d(n7953), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1710]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5882 (.d(n7954), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1709]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5883 (.d(n7955), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1708]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5884 (.d(n7956), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1707]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5885 (.d(n7957), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1706]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5886 (.d(n7958), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1705]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5887 (.d(n7959), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1704]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5888 (.d(n7960), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1703]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5889 (.d(n7961), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1702]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5890 (.d(n7962), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1701]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5891 (.d(n7963), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1700]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5892 (.d(n7964), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1699]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5893 (.d(n7965), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1698]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5894 (.d(n7966), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1697]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5895 (.d(n7967), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1696]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5896 (.d(n7968), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1695]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5897 (.d(n7969), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1694]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5898 (.d(n7970), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1693]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5899 (.d(n7971), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1692]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5900 (.d(n7972), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1691]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5901 (.d(n7973), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1690]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5902 (.d(n7974), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1689]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5903 (.d(n7975), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1688]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5904 (.d(n7976), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1687]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5905 (.d(n7977), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1686]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5906 (.d(n7978), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1685]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5907 (.d(n7979), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1684]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5908 (.d(n7980), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1683]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5909 (.d(n7981), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1682]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5910 (.d(n7982), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1681]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5911 (.d(n7983), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1680]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5912 (.d(n7984), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1679]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5913 (.d(n7985), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1678]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5914 (.d(n7986), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1677]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5915 (.d(n7987), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1676]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5916 (.d(n7988), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1675]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5917 (.d(n7989), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1674]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5918 (.d(n7990), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1673]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5919 (.d(n7991), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1672]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5920 (.d(n7992), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1671]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5921 (.d(n7993), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1670]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5922 (.d(n7994), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1669]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5923 (.d(n7995), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1668]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5924 (.d(n7996), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1667]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5925 (.d(n7997), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1666]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5926 (.d(n7998), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1665]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5927 (.d(n7999), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1664]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5928 (.d(n8000), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1663]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5929 (.d(n8001), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1662]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5930 (.d(n8002), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1661]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5931 (.d(n8003), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1660]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5932 (.d(n8004), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1659]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5933 (.d(n8005), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1658]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5934 (.d(n8006), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1657]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5935 (.d(n8007), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1656]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5936 (.d(n8008), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1655]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5937 (.d(n8009), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1654]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5938 (.d(n8010), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1653]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5939 (.d(n8011), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1652]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5940 (.d(n8012), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1651]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5941 (.d(n8013), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1650]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5942 (.d(n8014), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1649]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5943 (.d(n8015), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1648]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5944 (.d(n8016), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1647]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5945 (.d(n8017), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1646]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5946 (.d(n8018), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1645]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5947 (.d(n8019), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1644]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5948 (.d(n8020), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1643]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5949 (.d(n8021), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1642]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5950 (.d(n8022), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1641]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5951 (.d(n8023), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1640]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5952 (.d(n8024), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1639]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5953 (.d(n8025), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1638]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5954 (.d(n8026), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1637]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5955 (.d(n8027), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1636]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5956 (.d(n8028), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1635]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5957 (.d(n8029), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1634]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5958 (.d(n8030), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1633]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5959 (.d(n8031), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1632]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5960 (.d(n8032), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1631]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5961 (.d(n8033), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1630]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5962 (.d(n8034), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1629]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5963 (.d(n8035), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1628]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5964 (.d(n8036), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1627]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5965 (.d(n8037), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1626]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5966 (.d(n8038), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1625]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5967 (.d(n8039), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1624]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5968 (.d(n8040), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1623]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5969 (.d(n8041), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1622]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5970 (.d(n8042), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1621]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5971 (.d(n8043), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1620]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5972 (.d(n8044), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1619]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5973 (.d(n8045), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1618]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5974 (.d(n8046), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1617]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5975 (.d(n8047), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1616]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5976 (.d(n8048), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1615]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5977 (.d(n8049), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1614]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5978 (.d(n8050), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1613]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5979 (.d(n8051), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1612]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5980 (.d(n8052), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1611]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5981 (.d(n8053), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1610]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5982 (.d(n8054), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1609]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5983 (.d(n8055), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1608]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5984 (.d(n8056), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1607]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5985 (.d(n8057), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1606]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5986 (.d(n8058), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1605]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5987 (.d(n8059), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1604]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5988 (.d(n8060), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1603]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5989 (.d(n8061), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1602]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5990 (.d(n8062), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1601]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5991 (.d(n8063), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1600]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5992 (.d(n8064), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1599]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5993 (.d(n8065), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1598]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5994 (.d(n8066), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1597]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5995 (.d(n8067), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1596]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5996 (.d(n8068), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1595]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5997 (.d(n8069), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1594]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5998 (.d(n8070), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1593]));   // modexp_top.v(751)
    VERIFIC_DFFRS i5999 (.d(n8071), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1592]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6000 (.d(n8072), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1591]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6001 (.d(n8073), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1590]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6002 (.d(n8074), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1589]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6003 (.d(n8075), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1588]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6004 (.d(n8076), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1587]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6005 (.d(n8077), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1586]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6006 (.d(n8078), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1585]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6007 (.d(n8079), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1584]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6008 (.d(n8080), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1583]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6009 (.d(n8081), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1582]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6010 (.d(n8082), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1581]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6011 (.d(n8083), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1580]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6012 (.d(n8084), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1579]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6013 (.d(n8085), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1578]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6014 (.d(n8086), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1577]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6015 (.d(n8087), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1576]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6016 (.d(n8088), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1575]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6017 (.d(n8089), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1574]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6018 (.d(n8090), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1573]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6019 (.d(n8091), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1572]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6020 (.d(n8092), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1571]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6021 (.d(n8093), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1570]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6022 (.d(n8094), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1569]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6023 (.d(n8095), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1568]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6024 (.d(n8096), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1567]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6025 (.d(n8097), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1566]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6026 (.d(n8098), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1565]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6027 (.d(n8099), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1564]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6028 (.d(n8100), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1563]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6029 (.d(n8101), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1562]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6030 (.d(n8102), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1561]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6031 (.d(n8103), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1560]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6032 (.d(n8104), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1559]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6033 (.d(n8105), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1558]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6034 (.d(n8106), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1557]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6035 (.d(n8107), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1556]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6036 (.d(n8108), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1555]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6037 (.d(n8109), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1554]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6038 (.d(n8110), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1553]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6039 (.d(n8111), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1552]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6040 (.d(n8112), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1551]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6041 (.d(n8113), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1550]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6042 (.d(n8114), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1549]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6043 (.d(n8115), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1548]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6044 (.d(n8116), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1547]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6045 (.d(n8117), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1546]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6046 (.d(n8118), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1545]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6047 (.d(n8119), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1544]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6048 (.d(n8120), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1543]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6049 (.d(n8121), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1542]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6050 (.d(n8122), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1541]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6051 (.d(n8123), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1540]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6052 (.d(n8124), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1539]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6053 (.d(n8125), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1538]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6054 (.d(n8126), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1537]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6055 (.d(n8127), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1536]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6056 (.d(n8128), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1535]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6057 (.d(n8129), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1534]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6058 (.d(n8130), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1533]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6059 (.d(n8131), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1532]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6060 (.d(n8132), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1531]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6061 (.d(n8133), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1530]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6062 (.d(n8134), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1529]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6063 (.d(n8135), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1528]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6064 (.d(n8136), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1527]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6065 (.d(n8137), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1526]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6066 (.d(n8138), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1525]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6067 (.d(n8139), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1524]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6068 (.d(n8140), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1523]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6069 (.d(n8141), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1522]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6070 (.d(n8142), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1521]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6071 (.d(n8143), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1520]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6072 (.d(n8144), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1519]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6073 (.d(n8145), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1518]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6074 (.d(n8146), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1517]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6075 (.d(n8147), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1516]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6076 (.d(n8148), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1515]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6077 (.d(n8149), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1514]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6078 (.d(n8150), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1513]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6079 (.d(n8151), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1512]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6080 (.d(n8152), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1511]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6081 (.d(n8153), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1510]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6082 (.d(n8154), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1509]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6083 (.d(n8155), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1508]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6084 (.d(n8156), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1507]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6085 (.d(n8157), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1506]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6086 (.d(n8158), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1505]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6087 (.d(n8159), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1504]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6088 (.d(n8160), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1503]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6089 (.d(n8161), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1502]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6090 (.d(n8162), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1501]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6091 (.d(n8163), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1500]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6092 (.d(n8164), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1499]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6093 (.d(n8165), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1498]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6094 (.d(n8166), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1497]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6095 (.d(n8167), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1496]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6096 (.d(n8168), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1495]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6097 (.d(n8169), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1494]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6098 (.d(n8170), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1493]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6099 (.d(n8171), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1492]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6100 (.d(n8172), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1491]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6101 (.d(n8173), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1490]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6102 (.d(n8174), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1489]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6103 (.d(n8175), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1488]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6104 (.d(n8176), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1487]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6105 (.d(n8177), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1486]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6106 (.d(n8178), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1485]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6107 (.d(n8179), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1484]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6108 (.d(n8180), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1483]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6109 (.d(n8181), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1482]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6110 (.d(n8182), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1481]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6111 (.d(n8183), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1480]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6112 (.d(n8184), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1479]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6113 (.d(n8185), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1478]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6114 (.d(n8186), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1477]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6115 (.d(n8187), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1476]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6116 (.d(n8188), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1475]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6117 (.d(n8189), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1474]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6118 (.d(n8190), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1473]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6119 (.d(n8191), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1472]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6120 (.d(n8192), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1471]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6121 (.d(n8193), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1470]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6122 (.d(n8194), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1469]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6123 (.d(n8195), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1468]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6124 (.d(n8196), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1467]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6125 (.d(n8197), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1466]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6126 (.d(n8198), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1465]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6127 (.d(n8199), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1464]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6128 (.d(n8200), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1463]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6129 (.d(n8201), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1462]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6130 (.d(n8202), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1461]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6131 (.d(n8203), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1460]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6132 (.d(n8204), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1459]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6133 (.d(n8205), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1458]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6134 (.d(n8206), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1457]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6135 (.d(n8207), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1456]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6136 (.d(n8208), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1455]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6137 (.d(n8209), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1454]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6138 (.d(n8210), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1453]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6139 (.d(n8211), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1452]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6140 (.d(n8212), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1451]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6141 (.d(n8213), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1450]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6142 (.d(n8214), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1449]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6143 (.d(n8215), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1448]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6144 (.d(n8216), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1447]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6145 (.d(n8217), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1446]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6146 (.d(n8218), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1445]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6147 (.d(n8219), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1444]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6148 (.d(n8220), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1443]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6149 (.d(n8221), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1442]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6150 (.d(n8222), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1441]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6151 (.d(n8223), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1440]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6152 (.d(n8224), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1439]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6153 (.d(n8225), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1438]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6154 (.d(n8226), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1437]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6155 (.d(n8227), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1436]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6156 (.d(n8228), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1435]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6157 (.d(n8229), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1434]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6158 (.d(n8230), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1433]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6159 (.d(n8231), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1432]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6160 (.d(n8232), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1431]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6161 (.d(n8233), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1430]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6162 (.d(n8234), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1429]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6163 (.d(n8235), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1428]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6164 (.d(n8236), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1427]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6165 (.d(n8237), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1426]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6166 (.d(n8238), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1425]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6167 (.d(n8239), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1424]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6168 (.d(n8240), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1423]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6169 (.d(n8241), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1422]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6170 (.d(n8242), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1421]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6171 (.d(n8243), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1420]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6172 (.d(n8244), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1419]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6173 (.d(n8245), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1418]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6174 (.d(n8246), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1417]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6175 (.d(n8247), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1416]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6176 (.d(n8248), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1415]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6177 (.d(n8249), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1414]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6178 (.d(n8250), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1413]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6179 (.d(n8251), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1412]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6180 (.d(n8252), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1411]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6181 (.d(n8253), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1410]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6182 (.d(n8254), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1409]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6183 (.d(n8255), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1408]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6184 (.d(n8256), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1407]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6185 (.d(n8257), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1406]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6186 (.d(n8258), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1405]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6187 (.d(n8259), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1404]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6188 (.d(n8260), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1403]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6189 (.d(n8261), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1402]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6190 (.d(n8262), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1401]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6191 (.d(n8263), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1400]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6192 (.d(n8264), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1399]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6193 (.d(n8265), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1398]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6194 (.d(n8266), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1397]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6195 (.d(n8267), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1396]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6196 (.d(n8268), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1395]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6197 (.d(n8269), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1394]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6198 (.d(n8270), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1393]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6199 (.d(n8271), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1392]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6200 (.d(n8272), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1391]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6201 (.d(n8273), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1390]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6202 (.d(n8274), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1389]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6203 (.d(n8275), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1388]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6204 (.d(n8276), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1387]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6205 (.d(n8277), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1386]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6206 (.d(n8278), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1385]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6207 (.d(n8279), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1384]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6208 (.d(n8280), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1383]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6209 (.d(n8281), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1382]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6210 (.d(n8282), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1381]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6211 (.d(n8283), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1380]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6212 (.d(n8284), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1379]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6213 (.d(n8285), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1378]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6214 (.d(n8286), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1377]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6215 (.d(n8287), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1376]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6216 (.d(n8288), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1375]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6217 (.d(n8289), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1374]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6218 (.d(n8290), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1373]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6219 (.d(n8291), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1372]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6220 (.d(n8292), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1371]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6221 (.d(n8293), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1370]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6222 (.d(n8294), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1369]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6223 (.d(n8295), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1368]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6224 (.d(n8296), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1367]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6225 (.d(n8297), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1366]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6226 (.d(n8298), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1365]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6227 (.d(n8299), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1364]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6228 (.d(n8300), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1363]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6229 (.d(n8301), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1362]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6230 (.d(n8302), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1361]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6231 (.d(n8303), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1360]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6232 (.d(n8304), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1359]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6233 (.d(n8305), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1358]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6234 (.d(n8306), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1357]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6235 (.d(n8307), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1356]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6236 (.d(n8308), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1355]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6237 (.d(n8309), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1354]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6238 (.d(n8310), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1353]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6239 (.d(n8311), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1352]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6240 (.d(n8312), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1351]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6241 (.d(n8313), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1350]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6242 (.d(n8314), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1349]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6243 (.d(n8315), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1348]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6244 (.d(n8316), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1347]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6245 (.d(n8317), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1346]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6246 (.d(n8318), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1345]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6247 (.d(n8319), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1344]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6248 (.d(n8320), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1343]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6249 (.d(n8321), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1342]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6250 (.d(n8322), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1341]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6251 (.d(n8323), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1340]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6252 (.d(n8324), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1339]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6253 (.d(n8325), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1338]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6254 (.d(n8326), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1337]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6255 (.d(n8327), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1336]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6256 (.d(n8328), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1335]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6257 (.d(n8329), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1334]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6258 (.d(n8330), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1333]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6259 (.d(n8331), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1332]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6260 (.d(n8332), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1331]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6261 (.d(n8333), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1330]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6262 (.d(n8334), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1329]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6263 (.d(n8335), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1328]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6264 (.d(n8336), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1327]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6265 (.d(n8337), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1326]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6266 (.d(n8338), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1325]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6267 (.d(n8339), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1324]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6268 (.d(n8340), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1323]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6269 (.d(n8341), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1322]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6270 (.d(n8342), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1321]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6271 (.d(n8343), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1320]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6272 (.d(n8344), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1319]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6273 (.d(n8345), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1318]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6274 (.d(n8346), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1317]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6275 (.d(n8347), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1316]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6276 (.d(n8348), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1315]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6277 (.d(n8349), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1314]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6278 (.d(n8350), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1313]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6279 (.d(n8351), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1312]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6280 (.d(n8352), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1311]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6281 (.d(n8353), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1310]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6282 (.d(n8354), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1309]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6283 (.d(n8355), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1308]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6284 (.d(n8356), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1307]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6285 (.d(n8357), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1306]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6286 (.d(n8358), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1305]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6287 (.d(n8359), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1304]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6288 (.d(n8360), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1303]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6289 (.d(n8361), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1302]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6290 (.d(n8362), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1301]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6291 (.d(n8363), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1300]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6292 (.d(n8364), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1299]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6293 (.d(n8365), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1298]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6294 (.d(n8366), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1297]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6295 (.d(n8367), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1296]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6296 (.d(n8368), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1295]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6297 (.d(n8369), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1294]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6298 (.d(n8370), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1293]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6299 (.d(n8371), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1292]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6300 (.d(n8372), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1291]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6301 (.d(n8373), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1290]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6302 (.d(n8374), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1289]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6303 (.d(n8375), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1288]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6304 (.d(n8376), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1287]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6305 (.d(n8377), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1286]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6306 (.d(n8378), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1285]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6307 (.d(n8379), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1284]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6308 (.d(n8380), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1283]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6309 (.d(n8381), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1282]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6310 (.d(n8382), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1281]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6311 (.d(n8383), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1280]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6312 (.d(n8384), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1279]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6313 (.d(n8385), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1278]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6314 (.d(n8386), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1277]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6315 (.d(n8387), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1276]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6316 (.d(n8388), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1275]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6317 (.d(n8389), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1274]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6318 (.d(n8390), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1273]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6319 (.d(n8391), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1272]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6320 (.d(n8392), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1271]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6321 (.d(n8393), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1270]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6322 (.d(n8394), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1269]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6323 (.d(n8395), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1268]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6324 (.d(n8396), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1267]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6325 (.d(n8397), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1266]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6326 (.d(n8398), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1265]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6327 (.d(n8399), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1264]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6328 (.d(n8400), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1263]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6329 (.d(n8401), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1262]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6330 (.d(n8402), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1261]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6331 (.d(n8403), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1260]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6332 (.d(n8404), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1259]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6333 (.d(n8405), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1258]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6334 (.d(n8406), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1257]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6335 (.d(n8407), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1256]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6336 (.d(n8408), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1255]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6337 (.d(n8409), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1254]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6338 (.d(n8410), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1253]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6339 (.d(n8411), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1252]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6340 (.d(n8412), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1251]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6341 (.d(n8413), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1250]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6342 (.d(n8414), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1249]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6343 (.d(n8415), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1248]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6344 (.d(n8416), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1247]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6345 (.d(n8417), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1246]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6346 (.d(n8418), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1245]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6347 (.d(n8419), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1244]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6348 (.d(n8420), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1243]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6349 (.d(n8421), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1242]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6350 (.d(n8422), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1241]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6351 (.d(n8423), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1240]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6352 (.d(n8424), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1239]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6353 (.d(n8425), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1238]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6354 (.d(n8426), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1237]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6355 (.d(n8427), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1236]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6356 (.d(n8428), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1235]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6357 (.d(n8429), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1234]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6358 (.d(n8430), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1233]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6359 (.d(n8431), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1232]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6360 (.d(n8432), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1231]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6361 (.d(n8433), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1230]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6362 (.d(n8434), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1229]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6363 (.d(n8435), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1228]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6364 (.d(n8436), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1227]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6365 (.d(n8437), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1226]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6366 (.d(n8438), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1225]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6367 (.d(n8439), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1224]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6368 (.d(n8440), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1223]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6369 (.d(n8441), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1222]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6370 (.d(n8442), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1221]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6371 (.d(n8443), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1220]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6372 (.d(n8444), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1219]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6373 (.d(n8445), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1218]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6374 (.d(n8446), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1217]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6375 (.d(n8447), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1216]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6376 (.d(n8448), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1215]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6377 (.d(n8449), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1214]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6378 (.d(n8450), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1213]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6379 (.d(n8451), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1212]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6380 (.d(n8452), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1211]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6381 (.d(n8453), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1210]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6382 (.d(n8454), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1209]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6383 (.d(n8455), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1208]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6384 (.d(n8456), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1207]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6385 (.d(n8457), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1206]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6386 (.d(n8458), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1205]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6387 (.d(n8459), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1204]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6388 (.d(n8460), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1203]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6389 (.d(n8461), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1202]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6390 (.d(n8462), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1201]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6391 (.d(n8463), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1200]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6392 (.d(n8464), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1199]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6393 (.d(n8465), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1198]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6394 (.d(n8466), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1197]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6395 (.d(n8467), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1196]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6396 (.d(n8468), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1195]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6397 (.d(n8469), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1194]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6398 (.d(n8470), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1193]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6399 (.d(n8471), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1192]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6400 (.d(n8472), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1191]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6401 (.d(n8473), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1190]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6402 (.d(n8474), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1189]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6403 (.d(n8475), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1188]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6404 (.d(n8476), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1187]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6405 (.d(n8477), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1186]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6406 (.d(n8478), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1185]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6407 (.d(n8479), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1184]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6408 (.d(n8480), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1183]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6409 (.d(n8481), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1182]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6410 (.d(n8482), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1181]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6411 (.d(n8483), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1180]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6412 (.d(n8484), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1179]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6413 (.d(n8485), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1178]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6414 (.d(n8486), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1177]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6415 (.d(n8487), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1176]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6416 (.d(n8488), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1175]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6417 (.d(n8489), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1174]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6418 (.d(n8490), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1173]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6419 (.d(n8491), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1172]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6420 (.d(n8492), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1171]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6421 (.d(n8493), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1170]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6422 (.d(n8494), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1169]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6423 (.d(n8495), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1168]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6424 (.d(n8496), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1167]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6425 (.d(n8497), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1166]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6426 (.d(n8498), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1165]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6427 (.d(n8499), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1164]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6428 (.d(n8500), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1163]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6429 (.d(n8501), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1162]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6430 (.d(n8502), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1161]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6431 (.d(n8503), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1160]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6432 (.d(n8504), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1159]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6433 (.d(n8505), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1158]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6434 (.d(n8506), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1157]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6435 (.d(n8507), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1156]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6436 (.d(n8508), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1155]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6437 (.d(n8509), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1154]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6438 (.d(n8510), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1153]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6439 (.d(n8511), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1152]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6440 (.d(n8512), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1151]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6441 (.d(n8513), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1150]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6442 (.d(n8514), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1149]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6443 (.d(n8515), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1148]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6444 (.d(n8516), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1147]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6445 (.d(n8517), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1146]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6446 (.d(n8518), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1145]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6447 (.d(n8519), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1144]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6448 (.d(n8520), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1143]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6449 (.d(n8521), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1142]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6450 (.d(n8522), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1141]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6451 (.d(n8523), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1140]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6452 (.d(n8524), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1139]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6453 (.d(n8525), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1138]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6454 (.d(n8526), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1137]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6455 (.d(n8527), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1136]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6456 (.d(n8528), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1135]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6457 (.d(n8529), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1134]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6458 (.d(n8530), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1133]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6459 (.d(n8531), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1132]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6460 (.d(n8532), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1131]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6461 (.d(n8533), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1130]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6462 (.d(n8534), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1129]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6463 (.d(n8535), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1128]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6464 (.d(n8536), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1127]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6465 (.d(n8537), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1126]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6466 (.d(n8538), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1125]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6467 (.d(n8539), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1124]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6468 (.d(n8540), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1123]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6469 (.d(n8541), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1122]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6470 (.d(n8542), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1121]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6471 (.d(n8543), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1120]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6472 (.d(n8544), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1119]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6473 (.d(n8545), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1118]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6474 (.d(n8546), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1117]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6475 (.d(n8547), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1116]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6476 (.d(n8548), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1115]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6477 (.d(n8549), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1114]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6478 (.d(n8550), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1113]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6479 (.d(n8551), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1112]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6480 (.d(n8552), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1111]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6481 (.d(n8553), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1110]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6482 (.d(n8554), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1109]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6483 (.d(n8555), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1108]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6484 (.d(n8556), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1107]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6485 (.d(n8557), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1106]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6486 (.d(n8558), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1105]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6487 (.d(n8559), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1104]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6488 (.d(n8560), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1103]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6489 (.d(n8561), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1102]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6490 (.d(n8562), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1101]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6491 (.d(n8563), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1100]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6492 (.d(n8564), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1099]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6493 (.d(n8565), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1098]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6494 (.d(n8566), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1097]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6495 (.d(n8567), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1096]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6496 (.d(n8568), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1095]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6497 (.d(n8569), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1094]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6498 (.d(n8570), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1093]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6499 (.d(n8571), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1092]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6500 (.d(n8572), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1091]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6501 (.d(n8573), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1090]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6502 (.d(n8574), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1089]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6503 (.d(n8575), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1088]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6504 (.d(n8576), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1087]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6505 (.d(n8577), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1086]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6506 (.d(n8578), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1085]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6507 (.d(n8579), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1084]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6508 (.d(n8580), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1083]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6509 (.d(n8581), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1082]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6510 (.d(n8582), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1081]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6511 (.d(n8583), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1080]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6512 (.d(n8584), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1079]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6513 (.d(n8585), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1078]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6514 (.d(n8586), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1077]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6515 (.d(n8587), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1076]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6516 (.d(n8588), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1075]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6517 (.d(n8589), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1074]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6518 (.d(n8590), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1073]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6519 (.d(n8591), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1072]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6520 (.d(n8592), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1071]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6521 (.d(n8593), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1070]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6522 (.d(n8594), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1069]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6523 (.d(n8595), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1068]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6524 (.d(n8596), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1067]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6525 (.d(n8597), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1066]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6526 (.d(n8598), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1065]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6527 (.d(n8599), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1064]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6528 (.d(n8600), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1063]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6529 (.d(n8601), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1062]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6530 (.d(n8602), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1061]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6531 (.d(n8603), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1060]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6532 (.d(n8604), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1059]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6533 (.d(n8605), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1058]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6534 (.d(n8606), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1057]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6535 (.d(n8607), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1056]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6536 (.d(n8608), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1055]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6537 (.d(n8609), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1054]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6538 (.d(n8610), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1053]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6539 (.d(n8611), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1052]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6540 (.d(n8612), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1051]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6541 (.d(n8613), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1050]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6542 (.d(n8614), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1049]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6543 (.d(n8615), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1048]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6544 (.d(n8616), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1047]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6545 (.d(n8617), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1046]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6546 (.d(n8618), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1045]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6547 (.d(n8619), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1044]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6548 (.d(n8620), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1043]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6549 (.d(n8621), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1042]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6550 (.d(n8622), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1041]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6551 (.d(n8623), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1040]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6552 (.d(n8624), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1039]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6553 (.d(n8625), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1038]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6554 (.d(n8626), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1037]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6555 (.d(n8627), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1036]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6556 (.d(n8628), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1035]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6557 (.d(n8629), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1034]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6558 (.d(n8630), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1033]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6559 (.d(n8631), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1032]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6560 (.d(n8632), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1031]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6561 (.d(n8633), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1030]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6562 (.d(n8634), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1029]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6563 (.d(n8635), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1028]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6564 (.d(n8636), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1027]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6565 (.d(n8637), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1026]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6566 (.d(n8638), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1025]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6567 (.d(n8639), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1024]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6568 (.d(n8640), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1023]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6569 (.d(n8641), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1022]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6570 (.d(n8642), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1021]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6571 (.d(n8643), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1020]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6572 (.d(n8644), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1019]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6573 (.d(n8645), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1018]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6574 (.d(n8646), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1017]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6575 (.d(n8647), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1016]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6576 (.d(n8648), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1015]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6577 (.d(n8649), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1014]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6578 (.d(n8650), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1013]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6579 (.d(n8651), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1012]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6580 (.d(n8652), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1011]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6581 (.d(n8653), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1010]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6582 (.d(n8654), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1009]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6583 (.d(n8655), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1008]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6584 (.d(n8656), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1007]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6585 (.d(n8657), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1006]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6586 (.d(n8658), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1005]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6587 (.d(n8659), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1004]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6588 (.d(n8660), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1003]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6589 (.d(n8661), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1002]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6590 (.d(n8662), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1001]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6591 (.d(n8663), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1000]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6592 (.d(n8664), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[999]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6593 (.d(n8665), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[998]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6594 (.d(n8666), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[997]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6595 (.d(n8667), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[996]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6596 (.d(n8668), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[995]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6597 (.d(n8669), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[994]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6598 (.d(n8670), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[993]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6599 (.d(n8671), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[992]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6600 (.d(n8672), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[991]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6601 (.d(n8673), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[990]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6602 (.d(n8674), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[989]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6603 (.d(n8675), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[988]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6604 (.d(n8676), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[987]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6605 (.d(n8677), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[986]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6606 (.d(n8678), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[985]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6607 (.d(n8679), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[984]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6608 (.d(n8680), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[983]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6609 (.d(n8681), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[982]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6610 (.d(n8682), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[981]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6611 (.d(n8683), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[980]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6612 (.d(n8684), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[979]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6613 (.d(n8685), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[978]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6614 (.d(n8686), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[977]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6615 (.d(n8687), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[976]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6616 (.d(n8688), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[975]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6617 (.d(n8689), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[974]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6618 (.d(n8690), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[973]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6619 (.d(n8691), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[972]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6620 (.d(n8692), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[971]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6621 (.d(n8693), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[970]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6622 (.d(n8694), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[969]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6623 (.d(n8695), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[968]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6624 (.d(n8696), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[967]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6625 (.d(n8697), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[966]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6626 (.d(n8698), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[965]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6627 (.d(n8699), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[964]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6628 (.d(n8700), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[963]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6629 (.d(n8701), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[962]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6630 (.d(n8702), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[961]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6631 (.d(n8703), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[960]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6632 (.d(n8704), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[959]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6633 (.d(n8705), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[958]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6634 (.d(n8706), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[957]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6635 (.d(n8707), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[956]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6636 (.d(n8708), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[955]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6637 (.d(n8709), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[954]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6638 (.d(n8710), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[953]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6639 (.d(n8711), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[952]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6640 (.d(n8712), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[951]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6641 (.d(n8713), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[950]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6642 (.d(n8714), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[949]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6643 (.d(n8715), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[948]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6644 (.d(n8716), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[947]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6645 (.d(n8717), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[946]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6646 (.d(n8718), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[945]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6647 (.d(n8719), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[944]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6648 (.d(n8720), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[943]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6649 (.d(n8721), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[942]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6650 (.d(n8722), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[941]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6651 (.d(n8723), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[940]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6652 (.d(n8724), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[939]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6653 (.d(n8725), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[938]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6654 (.d(n8726), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[937]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6655 (.d(n8727), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[936]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6656 (.d(n8728), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[935]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6657 (.d(n8729), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[934]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6658 (.d(n8730), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[933]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6659 (.d(n8731), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[932]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6660 (.d(n8732), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[931]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6661 (.d(n8733), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[930]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6662 (.d(n8734), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[929]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6663 (.d(n8735), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[928]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6664 (.d(n8736), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[927]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6665 (.d(n8737), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[926]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6666 (.d(n8738), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[925]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6667 (.d(n8739), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[924]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6668 (.d(n8740), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[923]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6669 (.d(n8741), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[922]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6670 (.d(n8742), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[921]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6671 (.d(n8743), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[920]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6672 (.d(n8744), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[919]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6673 (.d(n8745), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[918]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6674 (.d(n8746), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[917]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6675 (.d(n8747), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[916]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6676 (.d(n8748), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[915]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6677 (.d(n8749), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[914]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6678 (.d(n8750), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[913]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6679 (.d(n8751), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[912]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6680 (.d(n8752), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[911]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6681 (.d(n8753), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[910]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6682 (.d(n8754), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[909]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6683 (.d(n8755), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[908]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6684 (.d(n8756), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[907]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6685 (.d(n8757), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[906]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6686 (.d(n8758), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[905]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6687 (.d(n8759), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[904]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6688 (.d(n8760), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[903]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6689 (.d(n8761), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[902]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6690 (.d(n8762), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[901]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6691 (.d(n8763), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[900]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6692 (.d(n8764), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[899]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6693 (.d(n8765), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[898]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6694 (.d(n8766), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[897]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6695 (.d(n8767), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[896]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6696 (.d(n8768), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[895]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6697 (.d(n8769), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[894]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6698 (.d(n8770), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[893]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6699 (.d(n8771), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[892]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6700 (.d(n8772), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[891]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6701 (.d(n8773), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[890]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6702 (.d(n8774), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[889]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6703 (.d(n8775), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[888]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6704 (.d(n8776), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[887]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6705 (.d(n8777), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[886]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6706 (.d(n8778), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[885]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6707 (.d(n8779), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[884]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6708 (.d(n8780), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[883]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6709 (.d(n8781), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[882]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6710 (.d(n8782), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[881]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6711 (.d(n8783), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[880]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6712 (.d(n8784), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[879]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6713 (.d(n8785), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[878]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6714 (.d(n8786), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[877]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6715 (.d(n8787), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[876]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6716 (.d(n8788), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[875]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6717 (.d(n8789), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[874]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6718 (.d(n8790), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[873]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6719 (.d(n8791), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[872]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6720 (.d(n8792), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[871]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6721 (.d(n8793), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[870]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6722 (.d(n8794), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[869]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6723 (.d(n8795), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[868]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6724 (.d(n8796), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[867]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6725 (.d(n8797), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[866]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6726 (.d(n8798), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[865]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6727 (.d(n8799), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[864]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6728 (.d(n8800), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[863]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6729 (.d(n8801), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[862]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6730 (.d(n8802), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[861]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6731 (.d(n8803), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[860]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6732 (.d(n8804), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[859]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6733 (.d(n8805), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[858]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6734 (.d(n8806), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[857]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6735 (.d(n8807), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[856]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6736 (.d(n8808), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[855]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6737 (.d(n8809), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[854]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6738 (.d(n8810), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[853]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6739 (.d(n8811), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[852]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6740 (.d(n8812), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[851]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6741 (.d(n8813), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[850]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6742 (.d(n8814), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[849]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6743 (.d(n8815), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[848]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6744 (.d(n8816), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[847]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6745 (.d(n8817), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[846]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6746 (.d(n8818), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[845]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6747 (.d(n8819), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[844]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6748 (.d(n8820), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[843]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6749 (.d(n8821), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[842]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6750 (.d(n8822), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[841]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6751 (.d(n8823), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[840]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6752 (.d(n8824), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[839]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6753 (.d(n8825), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[838]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6754 (.d(n8826), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[837]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6755 (.d(n8827), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[836]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6756 (.d(n8828), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[835]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6757 (.d(n8829), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[834]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6758 (.d(n8830), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[833]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6759 (.d(n8831), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[832]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6760 (.d(n8832), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[831]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6761 (.d(n8833), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[830]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6762 (.d(n8834), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[829]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6763 (.d(n8835), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[828]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6764 (.d(n8836), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[827]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6765 (.d(n8837), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[826]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6766 (.d(n8838), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[825]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6767 (.d(n8839), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[824]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6768 (.d(n8840), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[823]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6769 (.d(n8841), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[822]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6770 (.d(n8842), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[821]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6771 (.d(n8843), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[820]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6772 (.d(n8844), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[819]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6773 (.d(n8845), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[818]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6774 (.d(n8846), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[817]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6775 (.d(n8847), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[816]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6776 (.d(n8848), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[815]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6777 (.d(n8849), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[814]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6778 (.d(n8850), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[813]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6779 (.d(n8851), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[812]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6780 (.d(n8852), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[811]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6781 (.d(n8853), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[810]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6782 (.d(n8854), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[809]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6783 (.d(n8855), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[808]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6784 (.d(n8856), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[807]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6785 (.d(n8857), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[806]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6786 (.d(n8858), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[805]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6787 (.d(n8859), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[804]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6788 (.d(n8860), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[803]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6789 (.d(n8861), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[802]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6790 (.d(n8862), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[801]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6791 (.d(n8863), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[800]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6792 (.d(n8864), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[799]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6793 (.d(n8865), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[798]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6794 (.d(n8866), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[797]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6795 (.d(n8867), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[796]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6796 (.d(n8868), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[795]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6797 (.d(n8869), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[794]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6798 (.d(n8870), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[793]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6799 (.d(n8871), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[792]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6800 (.d(n8872), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[791]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6801 (.d(n8873), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[790]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6802 (.d(n8874), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[789]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6803 (.d(n8875), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[788]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6804 (.d(n8876), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[787]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6805 (.d(n8877), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[786]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6806 (.d(n8878), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[785]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6807 (.d(n8879), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[784]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6808 (.d(n8880), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[783]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6809 (.d(n8881), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[782]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6810 (.d(n8882), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[781]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6811 (.d(n8883), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[780]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6812 (.d(n8884), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[779]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6813 (.d(n8885), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[778]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6814 (.d(n8886), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[777]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6815 (.d(n8887), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[776]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6816 (.d(n8888), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[775]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6817 (.d(n8889), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[774]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6818 (.d(n8890), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[773]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6819 (.d(n8891), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[772]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6820 (.d(n8892), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[771]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6821 (.d(n8893), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[770]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6822 (.d(n8894), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[769]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6823 (.d(n8895), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[768]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6824 (.d(n8896), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[767]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6825 (.d(n8897), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[766]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6826 (.d(n8898), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[765]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6827 (.d(n8899), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[764]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6828 (.d(n8900), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[763]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6829 (.d(n8901), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[762]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6830 (.d(n8902), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[761]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6831 (.d(n8903), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[760]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6832 (.d(n8904), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[759]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6833 (.d(n8905), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[758]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6834 (.d(n8906), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[757]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6835 (.d(n8907), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[756]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6836 (.d(n8908), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[755]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6837 (.d(n8909), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[754]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6838 (.d(n8910), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[753]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6839 (.d(n8911), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[752]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6840 (.d(n8912), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[751]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6841 (.d(n8913), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[750]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6842 (.d(n8914), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[749]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6843 (.d(n8915), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[748]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6844 (.d(n8916), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[747]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6845 (.d(n8917), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[746]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6846 (.d(n8918), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[745]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6847 (.d(n8919), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[744]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6848 (.d(n8920), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[743]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6849 (.d(n8921), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[742]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6850 (.d(n8922), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[741]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6851 (.d(n8923), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[740]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6852 (.d(n8924), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[739]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6853 (.d(n8925), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[738]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6854 (.d(n8926), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[737]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6855 (.d(n8927), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[736]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6856 (.d(n8928), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[735]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6857 (.d(n8929), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[734]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6858 (.d(n8930), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[733]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6859 (.d(n8931), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[732]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6860 (.d(n8932), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[731]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6861 (.d(n8933), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[730]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6862 (.d(n8934), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[729]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6863 (.d(n8935), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[728]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6864 (.d(n8936), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[727]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6865 (.d(n8937), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[726]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6866 (.d(n8938), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[725]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6867 (.d(n8939), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[724]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6868 (.d(n8940), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[723]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6869 (.d(n8941), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[722]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6870 (.d(n8942), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[721]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6871 (.d(n8943), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[720]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6872 (.d(n8944), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[719]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6873 (.d(n8945), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[718]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6874 (.d(n8946), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[717]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6875 (.d(n8947), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[716]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6876 (.d(n8948), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[715]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6877 (.d(n8949), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[714]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6878 (.d(n8950), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[713]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6879 (.d(n8951), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[712]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6880 (.d(n8952), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[711]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6881 (.d(n8953), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[710]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6882 (.d(n8954), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[709]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6883 (.d(n8955), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[708]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6884 (.d(n8956), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[707]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6885 (.d(n8957), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[706]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6886 (.d(n8958), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[705]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6887 (.d(n8959), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[704]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6888 (.d(n8960), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[703]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6889 (.d(n8961), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[702]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6890 (.d(n8962), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[701]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6891 (.d(n8963), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[700]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6892 (.d(n8964), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[699]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6893 (.d(n8965), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[698]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6894 (.d(n8966), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[697]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6895 (.d(n8967), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[696]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6896 (.d(n8968), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[695]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6897 (.d(n8969), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[694]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6898 (.d(n8970), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[693]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6899 (.d(n8971), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[692]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6900 (.d(n8972), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[691]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6901 (.d(n8973), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[690]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6902 (.d(n8974), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[689]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6903 (.d(n8975), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[688]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6904 (.d(n8976), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[687]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6905 (.d(n8977), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[686]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6906 (.d(n8978), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[685]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6907 (.d(n8979), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[684]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6908 (.d(n8980), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[683]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6909 (.d(n8981), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[682]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6910 (.d(n8982), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[681]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6911 (.d(n8983), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[680]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6912 (.d(n8984), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[679]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6913 (.d(n8985), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[678]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6914 (.d(n8986), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[677]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6915 (.d(n8987), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[676]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6916 (.d(n8988), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[675]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6917 (.d(n8989), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[674]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6918 (.d(n8990), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[673]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6919 (.d(n8991), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[672]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6920 (.d(n8992), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[671]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6921 (.d(n8993), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[670]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6922 (.d(n8994), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[669]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6923 (.d(n8995), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[668]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6924 (.d(n8996), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[667]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6925 (.d(n8997), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[666]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6926 (.d(n8998), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[665]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6927 (.d(n8999), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[664]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6928 (.d(n9000), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[663]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6929 (.d(n9001), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[662]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6930 (.d(n9002), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[661]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6931 (.d(n9003), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[660]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6932 (.d(n9004), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[659]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6933 (.d(n9005), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[658]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6934 (.d(n9006), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[657]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6935 (.d(n9007), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[656]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6936 (.d(n9008), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[655]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6937 (.d(n9009), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[654]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6938 (.d(n9010), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[653]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6939 (.d(n9011), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[652]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6940 (.d(n9012), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[651]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6941 (.d(n9013), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[650]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6942 (.d(n9014), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[649]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6943 (.d(n9015), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[648]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6944 (.d(n9016), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[647]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6945 (.d(n9017), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[646]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6946 (.d(n9018), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[645]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6947 (.d(n9019), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[644]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6948 (.d(n9020), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[643]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6949 (.d(n9021), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[642]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6950 (.d(n9022), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[641]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6951 (.d(n9023), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[640]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6952 (.d(n9024), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[639]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6953 (.d(n9025), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[638]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6954 (.d(n9026), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[637]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6955 (.d(n9027), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[636]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6956 (.d(n9028), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[635]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6957 (.d(n9029), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[634]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6958 (.d(n9030), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[633]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6959 (.d(n9031), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[632]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6960 (.d(n9032), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[631]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6961 (.d(n9033), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[630]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6962 (.d(n9034), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[629]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6963 (.d(n9035), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[628]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6964 (.d(n9036), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[627]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6965 (.d(n9037), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[626]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6966 (.d(n9038), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[625]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6967 (.d(n9039), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[624]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6968 (.d(n9040), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[623]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6969 (.d(n9041), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[622]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6970 (.d(n9042), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[621]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6971 (.d(n9043), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[620]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6972 (.d(n9044), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[619]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6973 (.d(n9045), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[618]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6974 (.d(n9046), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[617]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6975 (.d(n9047), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[616]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6976 (.d(n9048), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[615]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6977 (.d(n9049), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[614]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6978 (.d(n9050), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[613]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6979 (.d(n9051), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[612]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6980 (.d(n9052), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[611]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6981 (.d(n9053), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[610]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6982 (.d(n9054), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[609]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6983 (.d(n9055), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[608]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6984 (.d(n9056), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[607]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6985 (.d(n9057), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[606]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6986 (.d(n9058), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[605]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6987 (.d(n9059), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[604]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6988 (.d(n9060), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[603]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6989 (.d(n9061), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[602]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6990 (.d(n9062), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[601]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6991 (.d(n9063), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[600]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6992 (.d(n9064), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[599]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6993 (.d(n9065), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[598]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6994 (.d(n9066), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[597]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6995 (.d(n9067), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[596]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6996 (.d(n9068), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[595]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6997 (.d(n9069), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[594]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6998 (.d(n9070), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[593]));   // modexp_top.v(751)
    VERIFIC_DFFRS i6999 (.d(n9071), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[592]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7000 (.d(n9072), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[591]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7001 (.d(n9073), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[590]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7002 (.d(n9074), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[589]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7003 (.d(n9075), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[588]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7004 (.d(n9076), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[587]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7005 (.d(n9077), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[586]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7006 (.d(n9078), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[585]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7007 (.d(n9079), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[584]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7008 (.d(n9080), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[583]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7009 (.d(n9081), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[582]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7010 (.d(n9082), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[581]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7011 (.d(n9083), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[580]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7012 (.d(n9084), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[579]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7013 (.d(n9085), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[578]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7014 (.d(n9086), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[577]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7015 (.d(n9087), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[576]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7016 (.d(n9088), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[575]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7017 (.d(n9089), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[574]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7018 (.d(n9090), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[573]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7019 (.d(n9091), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[572]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7020 (.d(n9092), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[571]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7021 (.d(n9093), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[570]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7022 (.d(n9094), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[569]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7023 (.d(n9095), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[568]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7024 (.d(n9096), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[567]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7025 (.d(n9097), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[566]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7026 (.d(n9098), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[565]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7027 (.d(n9099), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[564]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7028 (.d(n9100), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[563]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7029 (.d(n9101), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[562]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7030 (.d(n9102), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[561]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7031 (.d(n9103), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[560]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7032 (.d(n9104), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[559]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7033 (.d(n9105), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[558]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7034 (.d(n9106), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[557]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7035 (.d(n9107), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[556]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7036 (.d(n9108), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[555]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7037 (.d(n9109), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[554]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7038 (.d(n9110), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[553]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7039 (.d(n9111), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[552]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7040 (.d(n9112), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[551]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7041 (.d(n9113), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[550]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7042 (.d(n9114), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[549]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7043 (.d(n9115), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[548]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7044 (.d(n9116), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[547]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7045 (.d(n9117), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[546]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7046 (.d(n9118), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[545]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7047 (.d(n9119), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[544]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7048 (.d(n9120), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[543]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7049 (.d(n9121), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[542]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7050 (.d(n9122), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[541]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7051 (.d(n9123), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[540]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7052 (.d(n9124), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[539]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7053 (.d(n9125), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[538]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7054 (.d(n9126), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[537]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7055 (.d(n9127), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[536]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7056 (.d(n9128), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[535]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7057 (.d(n9129), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[534]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7058 (.d(n9130), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[533]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7059 (.d(n9131), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[532]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7060 (.d(n9132), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[531]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7061 (.d(n9133), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[530]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7062 (.d(n9134), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[529]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7063 (.d(n9135), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[528]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7064 (.d(n9136), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[527]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7065 (.d(n9137), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[526]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7066 (.d(n9138), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[525]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7067 (.d(n9139), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[524]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7068 (.d(n9140), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[523]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7069 (.d(n9141), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[522]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7070 (.d(n9142), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[521]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7071 (.d(n9143), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[520]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7072 (.d(n9144), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[519]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7073 (.d(n9145), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[518]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7074 (.d(n9146), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[517]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7075 (.d(n9147), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[516]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7076 (.d(n9148), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[515]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7077 (.d(n9149), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[514]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7078 (.d(n9150), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[513]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7079 (.d(n9151), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[512]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7080 (.d(n9152), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[511]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7081 (.d(n9153), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[510]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7082 (.d(n9154), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[509]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7083 (.d(n9155), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[508]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7084 (.d(n9156), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[507]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7085 (.d(n9157), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[506]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7086 (.d(n9158), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[505]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7087 (.d(n9159), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[504]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7088 (.d(n9160), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[503]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7089 (.d(n9161), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[502]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7090 (.d(n9162), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[501]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7091 (.d(n9163), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[500]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7092 (.d(n9164), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[499]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7093 (.d(n9165), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[498]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7094 (.d(n9166), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[497]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7095 (.d(n9167), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[496]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7096 (.d(n9168), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[495]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7097 (.d(n9169), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[494]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7098 (.d(n9170), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[493]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7099 (.d(n9171), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[492]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7100 (.d(n9172), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[491]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7101 (.d(n9173), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[490]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7102 (.d(n9174), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[489]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7103 (.d(n9175), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[488]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7104 (.d(n9176), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[487]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7105 (.d(n9177), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[486]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7106 (.d(n9178), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[485]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7107 (.d(n9179), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[484]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7108 (.d(n9180), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[483]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7109 (.d(n9181), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[482]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7110 (.d(n9182), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[481]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7111 (.d(n9183), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[480]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7112 (.d(n9184), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[479]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7113 (.d(n9185), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[478]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7114 (.d(n9186), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[477]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7115 (.d(n9187), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[476]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7116 (.d(n9188), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[475]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7117 (.d(n9189), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[474]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7118 (.d(n9190), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[473]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7119 (.d(n9191), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[472]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7120 (.d(n9192), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[471]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7121 (.d(n9193), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[470]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7122 (.d(n9194), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[469]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7123 (.d(n9195), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[468]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7124 (.d(n9196), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[467]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7125 (.d(n9197), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[466]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7126 (.d(n9198), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[465]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7127 (.d(n9199), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[464]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7128 (.d(n9200), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[463]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7129 (.d(n9201), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[462]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7130 (.d(n9202), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[461]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7131 (.d(n9203), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[460]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7132 (.d(n9204), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[459]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7133 (.d(n9205), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[458]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7134 (.d(n9206), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[457]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7135 (.d(n9207), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[456]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7136 (.d(n9208), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[455]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7137 (.d(n9209), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[454]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7138 (.d(n9210), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[453]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7139 (.d(n9211), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[452]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7140 (.d(n9212), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[451]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7141 (.d(n9213), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[450]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7142 (.d(n9214), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[449]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7143 (.d(n9215), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[448]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7144 (.d(n9216), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[447]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7145 (.d(n9217), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[446]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7146 (.d(n9218), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[445]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7147 (.d(n9219), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[444]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7148 (.d(n9220), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[443]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7149 (.d(n9221), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[442]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7150 (.d(n9222), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[441]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7151 (.d(n9223), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[440]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7152 (.d(n9224), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[439]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7153 (.d(n9225), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[438]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7154 (.d(n9226), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[437]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7155 (.d(n9227), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[436]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7156 (.d(n9228), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[435]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7157 (.d(n9229), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[434]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7158 (.d(n9230), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[433]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7159 (.d(n9231), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[432]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7160 (.d(n9232), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[431]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7161 (.d(n9233), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[430]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7162 (.d(n9234), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[429]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7163 (.d(n9235), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[428]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7164 (.d(n9236), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[427]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7165 (.d(n9237), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[426]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7166 (.d(n9238), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[425]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7167 (.d(n9239), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[424]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7168 (.d(n9240), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[423]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7169 (.d(n9241), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[422]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7170 (.d(n9242), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[421]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7171 (.d(n9243), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[420]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7172 (.d(n9244), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[419]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7173 (.d(n9245), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[418]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7174 (.d(n9246), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[417]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7175 (.d(n9247), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[416]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7176 (.d(n9248), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[415]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7177 (.d(n9249), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[414]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7178 (.d(n9250), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[413]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7179 (.d(n9251), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[412]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7180 (.d(n9252), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[411]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7181 (.d(n9253), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[410]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7182 (.d(n9254), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[409]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7183 (.d(n9255), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[408]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7184 (.d(n9256), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[407]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7185 (.d(n9257), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[406]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7186 (.d(n9258), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[405]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7187 (.d(n9259), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[404]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7188 (.d(n9260), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[403]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7189 (.d(n9261), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[402]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7190 (.d(n9262), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[401]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7191 (.d(n9263), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[400]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7192 (.d(n9264), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[399]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7193 (.d(n9265), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[398]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7194 (.d(n9266), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[397]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7195 (.d(n9267), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[396]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7196 (.d(n9268), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[395]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7197 (.d(n9269), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[394]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7198 (.d(n9270), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[393]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7199 (.d(n9271), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[392]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7200 (.d(n9272), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[391]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7201 (.d(n9273), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[390]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7202 (.d(n9274), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[389]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7203 (.d(n9275), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[388]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7204 (.d(n9276), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[387]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7205 (.d(n9277), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[386]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7206 (.d(n9278), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[385]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7207 (.d(n9279), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[384]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7208 (.d(n9280), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[383]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7209 (.d(n9281), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[382]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7210 (.d(n9282), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[381]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7211 (.d(n9283), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[380]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7212 (.d(n9284), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[379]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7213 (.d(n9285), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[378]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7214 (.d(n9286), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[377]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7215 (.d(n9287), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[376]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7216 (.d(n9288), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[375]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7217 (.d(n9289), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[374]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7218 (.d(n9290), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[373]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7219 (.d(n9291), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[372]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7220 (.d(n9292), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[371]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7221 (.d(n9293), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[370]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7222 (.d(n9294), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[369]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7223 (.d(n9295), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[368]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7224 (.d(n9296), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[367]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7225 (.d(n9297), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[366]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7226 (.d(n9298), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[365]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7227 (.d(n9299), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[364]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7228 (.d(n9300), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[363]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7229 (.d(n9301), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[362]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7230 (.d(n9302), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[361]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7231 (.d(n9303), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[360]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7232 (.d(n9304), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[359]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7233 (.d(n9305), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[358]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7234 (.d(n9306), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[357]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7235 (.d(n9307), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[356]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7236 (.d(n9308), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[355]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7237 (.d(n9309), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[354]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7238 (.d(n9310), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[353]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7239 (.d(n9311), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[352]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7240 (.d(n9312), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[351]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7241 (.d(n9313), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[350]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7242 (.d(n9314), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[349]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7243 (.d(n9315), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[348]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7244 (.d(n9316), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[347]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7245 (.d(n9317), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[346]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7246 (.d(n9318), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[345]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7247 (.d(n9319), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[344]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7248 (.d(n9320), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[343]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7249 (.d(n9321), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[342]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7250 (.d(n9322), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[341]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7251 (.d(n9323), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[340]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7252 (.d(n9324), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[339]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7253 (.d(n9325), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[338]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7254 (.d(n9326), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[337]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7255 (.d(n9327), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[336]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7256 (.d(n9328), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[335]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7257 (.d(n9329), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[334]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7258 (.d(n9330), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[333]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7259 (.d(n9331), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[332]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7260 (.d(n9332), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[331]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7261 (.d(n9333), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[330]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7262 (.d(n9334), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[329]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7263 (.d(n9335), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[328]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7264 (.d(n9336), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[327]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7265 (.d(n9337), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[326]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7266 (.d(n9338), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[325]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7267 (.d(n9339), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[324]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7268 (.d(n9340), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[323]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7269 (.d(n9341), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[322]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7270 (.d(n9342), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[321]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7271 (.d(n9343), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[320]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7272 (.d(n9344), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[319]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7273 (.d(n9345), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[318]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7274 (.d(n9346), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[317]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7275 (.d(n9347), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[316]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7276 (.d(n9348), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[315]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7277 (.d(n9349), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[314]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7278 (.d(n9350), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[313]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7279 (.d(n9351), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[312]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7280 (.d(n9352), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[311]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7281 (.d(n9353), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[310]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7282 (.d(n9354), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[309]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7283 (.d(n9355), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[308]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7284 (.d(n9356), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[307]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7285 (.d(n9357), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[306]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7286 (.d(n9358), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[305]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7287 (.d(n9359), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[304]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7288 (.d(n9360), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[303]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7289 (.d(n9361), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[302]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7290 (.d(n9362), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[301]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7291 (.d(n9363), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[300]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7292 (.d(n9364), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[299]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7293 (.d(n9365), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[298]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7294 (.d(n9366), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[297]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7295 (.d(n9367), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[296]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7296 (.d(n9368), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[295]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7297 (.d(n9369), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[294]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7298 (.d(n9370), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[293]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7299 (.d(n9371), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[292]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7300 (.d(n9372), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[291]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7301 (.d(n9373), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[290]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7302 (.d(n9374), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[289]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7303 (.d(n9375), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[288]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7304 (.d(n9376), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[287]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7305 (.d(n9377), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[286]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7306 (.d(n9378), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[285]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7307 (.d(n9379), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[284]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7308 (.d(n9380), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[283]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7309 (.d(n9381), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[282]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7310 (.d(n9382), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[281]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7311 (.d(n9383), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[280]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7312 (.d(n9384), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[279]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7313 (.d(n9385), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[278]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7314 (.d(n9386), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[277]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7315 (.d(n9387), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[276]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7316 (.d(n9388), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[275]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7317 (.d(n9389), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[274]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7318 (.d(n9390), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[273]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7319 (.d(n9391), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[272]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7320 (.d(n9392), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[271]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7321 (.d(n9393), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[270]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7322 (.d(n9394), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[269]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7323 (.d(n9395), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[268]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7324 (.d(n9396), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[267]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7325 (.d(n9397), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[266]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7326 (.d(n9398), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[265]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7327 (.d(n9399), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[264]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7328 (.d(n9400), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[263]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7329 (.d(n9401), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[262]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7330 (.d(n9402), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[261]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7331 (.d(n9403), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[260]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7332 (.d(n9404), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[259]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7333 (.d(n9405), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[258]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7334 (.d(n9406), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[257]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7335 (.d(n9407), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[256]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7336 (.d(n9408), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[255]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7337 (.d(n9409), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[254]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7338 (.d(n9410), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[253]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7339 (.d(n9411), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[252]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7340 (.d(n9412), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[251]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7341 (.d(n9413), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[250]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7342 (.d(n9414), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[249]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7343 (.d(n9415), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[248]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7344 (.d(n9416), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[247]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7345 (.d(n9417), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[246]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7346 (.d(n9418), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[245]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7347 (.d(n9419), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[244]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7348 (.d(n9420), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[243]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7349 (.d(n9421), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[242]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7350 (.d(n9422), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[241]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7351 (.d(n9423), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[240]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7352 (.d(n9424), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[239]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7353 (.d(n9425), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[238]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7354 (.d(n9426), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[237]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7355 (.d(n9427), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[236]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7356 (.d(n9428), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[235]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7357 (.d(n9429), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[234]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7358 (.d(n9430), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[233]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7359 (.d(n9431), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[232]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7360 (.d(n9432), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[231]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7361 (.d(n9433), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[230]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7362 (.d(n9434), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[229]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7363 (.d(n9435), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[228]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7364 (.d(n9436), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[227]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7365 (.d(n9437), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[226]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7366 (.d(n9438), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[225]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7367 (.d(n9439), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[224]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7368 (.d(n9440), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[223]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7369 (.d(n9441), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[222]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7370 (.d(n9442), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[221]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7371 (.d(n9443), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[220]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7372 (.d(n9444), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[219]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7373 (.d(n9445), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[218]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7374 (.d(n9446), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[217]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7375 (.d(n9447), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[216]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7376 (.d(n9448), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[215]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7377 (.d(n9449), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[214]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7378 (.d(n9450), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[213]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7379 (.d(n9451), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[212]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7380 (.d(n9452), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[211]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7381 (.d(n9453), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[210]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7382 (.d(n9454), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[209]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7383 (.d(n9455), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[208]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7384 (.d(n9456), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[207]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7385 (.d(n9457), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[206]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7386 (.d(n9458), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[205]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7387 (.d(n9459), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[204]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7388 (.d(n9460), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[203]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7389 (.d(n9461), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[202]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7390 (.d(n9462), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[201]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7391 (.d(n9463), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[200]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7392 (.d(n9464), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[199]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7393 (.d(n9465), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[198]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7394 (.d(n9466), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[197]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7395 (.d(n9467), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[196]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7396 (.d(n9468), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[195]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7397 (.d(n9469), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[194]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7398 (.d(n9470), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[193]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7399 (.d(n9471), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[192]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7400 (.d(n9472), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[191]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7401 (.d(n9473), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[190]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7402 (.d(n9474), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[189]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7403 (.d(n9475), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[188]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7404 (.d(n9476), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[187]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7405 (.d(n9477), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[186]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7406 (.d(n9478), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[185]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7407 (.d(n9479), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[184]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7408 (.d(n9480), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[183]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7409 (.d(n9481), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[182]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7410 (.d(n9482), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[181]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7411 (.d(n9483), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[180]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7412 (.d(n9484), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[179]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7413 (.d(n9485), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[178]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7414 (.d(n9486), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[177]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7415 (.d(n9487), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[176]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7416 (.d(n9488), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[175]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7417 (.d(n9489), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[174]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7418 (.d(n9490), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[173]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7419 (.d(n9491), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[172]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7420 (.d(n9492), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[171]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7421 (.d(n9493), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[170]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7422 (.d(n9494), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[169]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7423 (.d(n9495), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[168]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7424 (.d(n9496), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[167]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7425 (.d(n9497), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[166]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7426 (.d(n9498), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[165]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7427 (.d(n9499), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[164]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7428 (.d(n9500), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[163]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7429 (.d(n9501), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[162]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7430 (.d(n9502), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[161]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7431 (.d(n9503), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[160]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7432 (.d(n9504), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[159]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7433 (.d(n9505), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[158]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7434 (.d(n9506), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[157]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7435 (.d(n9507), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[156]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7436 (.d(n9508), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[155]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7437 (.d(n9509), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[154]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7438 (.d(n9510), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[153]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7439 (.d(n9511), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[152]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7440 (.d(n9512), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[151]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7441 (.d(n9513), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[150]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7442 (.d(n9514), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[149]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7443 (.d(n9515), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[148]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7444 (.d(n9516), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[147]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7445 (.d(n9517), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[146]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7446 (.d(n9518), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[145]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7447 (.d(n9519), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[144]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7448 (.d(n9520), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[143]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7449 (.d(n9521), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[142]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7450 (.d(n9522), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[141]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7451 (.d(n9523), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[140]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7452 (.d(n9524), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[139]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7453 (.d(n9525), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[138]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7454 (.d(n9526), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[137]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7455 (.d(n9527), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[136]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7456 (.d(n9528), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[135]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7457 (.d(n9529), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[134]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7458 (.d(n9530), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[133]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7459 (.d(n9531), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[132]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7460 (.d(n9532), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[131]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7461 (.d(n9533), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[130]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7462 (.d(n9534), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[129]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7463 (.d(n9535), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[128]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7464 (.d(n9536), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[127]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7465 (.d(n9537), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[126]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7466 (.d(n9538), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[125]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7467 (.d(n9539), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[124]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7468 (.d(n9540), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[123]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7469 (.d(n9541), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[122]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7470 (.d(n9542), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[121]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7471 (.d(n9543), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[120]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7472 (.d(n9544), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[119]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7473 (.d(n9545), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[118]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7474 (.d(n9546), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[117]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7475 (.d(n9547), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[116]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7476 (.d(n9548), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[115]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7477 (.d(n9549), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[114]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7478 (.d(n9550), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[113]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7479 (.d(n9551), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[112]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7480 (.d(n9552), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[111]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7481 (.d(n9553), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[110]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7482 (.d(n9554), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[109]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7483 (.d(n9555), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[108]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7484 (.d(n9556), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[107]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7485 (.d(n9557), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[106]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7486 (.d(n9558), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[105]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7487 (.d(n9559), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[104]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7488 (.d(n9560), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[103]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7489 (.d(n9561), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[102]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7490 (.d(n9562), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[101]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7491 (.d(n9563), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[100]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7492 (.d(n9564), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[99]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7493 (.d(n9565), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[98]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7494 (.d(n9566), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[97]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7495 (.d(n9567), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[96]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7496 (.d(n9568), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[95]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7497 (.d(n9569), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[94]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7498 (.d(n9570), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[93]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7499 (.d(n9571), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[92]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7500 (.d(n9572), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[91]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7501 (.d(n9573), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[90]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7502 (.d(n9574), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[89]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7503 (.d(n9575), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[88]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7504 (.d(n9576), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[87]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7505 (.d(n9577), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[86]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7506 (.d(n9578), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[85]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7507 (.d(n9579), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[84]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7508 (.d(n9580), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[83]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7509 (.d(n9581), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[82]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7510 (.d(n9582), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[81]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7511 (.d(n9583), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[80]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7512 (.d(n9584), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[79]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7513 (.d(n9585), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[78]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7514 (.d(n9586), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[77]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7515 (.d(n9587), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[76]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7516 (.d(n9588), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[75]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7517 (.d(n9589), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[74]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7518 (.d(n9590), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[73]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7519 (.d(n9591), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[72]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7520 (.d(n9592), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[71]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7521 (.d(n9593), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[70]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7522 (.d(n9594), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[69]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7523 (.d(n9595), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[68]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7524 (.d(n9596), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[67]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7525 (.d(n9597), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[66]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7526 (.d(n9598), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[65]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7527 (.d(n9599), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[64]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7528 (.d(n9600), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[63]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7529 (.d(n9601), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[62]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7530 (.d(n9602), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[61]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7531 (.d(n9603), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[60]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7532 (.d(n9604), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[59]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7533 (.d(n9605), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[58]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7534 (.d(n9606), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[57]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7535 (.d(n9607), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[56]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7536 (.d(n9608), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[55]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7537 (.d(n9609), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[54]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7538 (.d(n9610), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[53]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7539 (.d(n9611), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[52]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7540 (.d(n9612), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[51]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7541 (.d(n9613), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[50]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7542 (.d(n9614), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[49]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7543 (.d(n9615), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[48]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7544 (.d(n9616), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[47]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7545 (.d(n9617), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[46]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7546 (.d(n9618), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[45]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7547 (.d(n9619), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[44]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7548 (.d(n9620), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[43]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7549 (.d(n9621), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[42]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7550 (.d(n9622), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[41]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7551 (.d(n9623), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[40]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7552 (.d(n9624), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[39]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7553 (.d(n9625), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[38]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7554 (.d(n9626), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[37]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7555 (.d(n9627), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[36]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7556 (.d(n9628), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[35]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7557 (.d(n9629), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[34]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7558 (.d(n9630), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[33]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7559 (.d(n9631), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[32]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7560 (.d(n9632), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[31]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7561 (.d(n9633), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[30]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7562 (.d(n9634), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[29]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7563 (.d(n9635), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[28]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7564 (.d(n9636), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[27]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7565 (.d(n9637), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[26]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7566 (.d(n9638), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[25]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7567 (.d(n9639), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[24]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7568 (.d(n9640), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[23]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7569 (.d(n9641), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[22]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7570 (.d(n9642), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[21]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7571 (.d(n9643), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[20]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7572 (.d(n9644), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[19]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7573 (.d(n9645), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[18]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7574 (.d(n9646), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[17]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7575 (.d(n9647), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[16]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7576 (.d(n9648), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[15]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7577 (.d(n9649), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[14]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7578 (.d(n9650), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[13]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7579 (.d(n9651), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[12]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7580 (.d(n9652), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[11]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7581 (.d(n9653), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[10]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7582 (.d(n9654), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[9]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7583 (.d(n9655), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[8]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7584 (.d(n9656), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[7]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7585 (.d(n9657), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[6]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7586 (.d(n9658), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[5]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7587 (.d(n9659), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[4]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7588 (.d(n9660), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[3]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7589 (.d(n9661), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[2]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7590 (.d(n9662), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[1]));   // modexp_top.v(751)
    VERIFIC_DFFRS i7591 (.d(n9663), .clk(clk), .s(1'b0), .r(1'b0), .q(encrypted_data_buf[0]));   // modexp_top.v(751)
    assign n7616 = rst ? encrypted_data_buf[2047] : encrypted_data_buf_next[2047];   // modexp_top.v(751)
    assign n7617 = rst ? encrypted_data_buf[2046] : encrypted_data_buf_next[2046];   // modexp_top.v(751)
    assign n7618 = rst ? encrypted_data_buf[2045] : encrypted_data_buf_next[2045];   // modexp_top.v(751)
    assign n7619 = rst ? encrypted_data_buf[2044] : encrypted_data_buf_next[2044];   // modexp_top.v(751)
    assign n7620 = rst ? encrypted_data_buf[2043] : encrypted_data_buf_next[2043];   // modexp_top.v(751)
    assign n7621 = rst ? encrypted_data_buf[2042] : encrypted_data_buf_next[2042];   // modexp_top.v(751)
    assign n7622 = rst ? encrypted_data_buf[2041] : encrypted_data_buf_next[2041];   // modexp_top.v(751)
    assign n7623 = rst ? encrypted_data_buf[2040] : encrypted_data_buf_next[2040];   // modexp_top.v(751)
    assign n7624 = rst ? encrypted_data_buf[2039] : encrypted_data_buf_next[2039];   // modexp_top.v(751)
    assign n7625 = rst ? encrypted_data_buf[2038] : encrypted_data_buf_next[2038];   // modexp_top.v(751)
    assign n7626 = rst ? encrypted_data_buf[2037] : encrypted_data_buf_next[2037];   // modexp_top.v(751)
    assign n7627 = rst ? encrypted_data_buf[2036] : encrypted_data_buf_next[2036];   // modexp_top.v(751)
    assign n7628 = rst ? encrypted_data_buf[2035] : encrypted_data_buf_next[2035];   // modexp_top.v(751)
    assign n7629 = rst ? encrypted_data_buf[2034] : encrypted_data_buf_next[2034];   // modexp_top.v(751)
    assign n7630 = rst ? encrypted_data_buf[2033] : encrypted_data_buf_next[2033];   // modexp_top.v(751)
    assign n7631 = rst ? encrypted_data_buf[2032] : encrypted_data_buf_next[2032];   // modexp_top.v(751)
    assign n7632 = rst ? encrypted_data_buf[2031] : encrypted_data_buf_next[2031];   // modexp_top.v(751)
    assign n7633 = rst ? encrypted_data_buf[2030] : encrypted_data_buf_next[2030];   // modexp_top.v(751)
    assign n7634 = rst ? encrypted_data_buf[2029] : encrypted_data_buf_next[2029];   // modexp_top.v(751)
    assign n7635 = rst ? encrypted_data_buf[2028] : encrypted_data_buf_next[2028];   // modexp_top.v(751)
    assign n7636 = rst ? encrypted_data_buf[2027] : encrypted_data_buf_next[2027];   // modexp_top.v(751)
    assign n7637 = rst ? encrypted_data_buf[2026] : encrypted_data_buf_next[2026];   // modexp_top.v(751)
    assign n7638 = rst ? encrypted_data_buf[2025] : encrypted_data_buf_next[2025];   // modexp_top.v(751)
    assign n7639 = rst ? encrypted_data_buf[2024] : encrypted_data_buf_next[2024];   // modexp_top.v(751)
    assign n7640 = rst ? encrypted_data_buf[2023] : encrypted_data_buf_next[2023];   // modexp_top.v(751)
    assign n7641 = rst ? encrypted_data_buf[2022] : encrypted_data_buf_next[2022];   // modexp_top.v(751)
    assign n7642 = rst ? encrypted_data_buf[2021] : encrypted_data_buf_next[2021];   // modexp_top.v(751)
    assign n7643 = rst ? encrypted_data_buf[2020] : encrypted_data_buf_next[2020];   // modexp_top.v(751)
    assign n7644 = rst ? encrypted_data_buf[2019] : encrypted_data_buf_next[2019];   // modexp_top.v(751)
    assign n7645 = rst ? encrypted_data_buf[2018] : encrypted_data_buf_next[2018];   // modexp_top.v(751)
    assign n7646 = rst ? encrypted_data_buf[2017] : encrypted_data_buf_next[2017];   // modexp_top.v(751)
    assign n7647 = rst ? encrypted_data_buf[2016] : encrypted_data_buf_next[2016];   // modexp_top.v(751)
    assign n7648 = rst ? encrypted_data_buf[2015] : encrypted_data_buf_next[2015];   // modexp_top.v(751)
    assign n7649 = rst ? encrypted_data_buf[2014] : encrypted_data_buf_next[2014];   // modexp_top.v(751)
    assign n7650 = rst ? encrypted_data_buf[2013] : encrypted_data_buf_next[2013];   // modexp_top.v(751)
    assign n7651 = rst ? encrypted_data_buf[2012] : encrypted_data_buf_next[2012];   // modexp_top.v(751)
    assign n7652 = rst ? encrypted_data_buf[2011] : encrypted_data_buf_next[2011];   // modexp_top.v(751)
    assign n7653 = rst ? encrypted_data_buf[2010] : encrypted_data_buf_next[2010];   // modexp_top.v(751)
    assign n7654 = rst ? encrypted_data_buf[2009] : encrypted_data_buf_next[2009];   // modexp_top.v(751)
    assign n7655 = rst ? encrypted_data_buf[2008] : encrypted_data_buf_next[2008];   // modexp_top.v(751)
    assign n7656 = rst ? encrypted_data_buf[2007] : encrypted_data_buf_next[2007];   // modexp_top.v(751)
    assign n7657 = rst ? encrypted_data_buf[2006] : encrypted_data_buf_next[2006];   // modexp_top.v(751)
    assign n7658 = rst ? encrypted_data_buf[2005] : encrypted_data_buf_next[2005];   // modexp_top.v(751)
    assign n7659 = rst ? encrypted_data_buf[2004] : encrypted_data_buf_next[2004];   // modexp_top.v(751)
    assign n7660 = rst ? encrypted_data_buf[2003] : encrypted_data_buf_next[2003];   // modexp_top.v(751)
    assign n7661 = rst ? encrypted_data_buf[2002] : encrypted_data_buf_next[2002];   // modexp_top.v(751)
    assign n7662 = rst ? encrypted_data_buf[2001] : encrypted_data_buf_next[2001];   // modexp_top.v(751)
    assign n7663 = rst ? encrypted_data_buf[2000] : encrypted_data_buf_next[2000];   // modexp_top.v(751)
    assign n7664 = rst ? encrypted_data_buf[1999] : encrypted_data_buf_next[1999];   // modexp_top.v(751)
    assign n7665 = rst ? encrypted_data_buf[1998] : encrypted_data_buf_next[1998];   // modexp_top.v(751)
    assign n7666 = rst ? encrypted_data_buf[1997] : encrypted_data_buf_next[1997];   // modexp_top.v(751)
    assign n7667 = rst ? encrypted_data_buf[1996] : encrypted_data_buf_next[1996];   // modexp_top.v(751)
    assign n7668 = rst ? encrypted_data_buf[1995] : encrypted_data_buf_next[1995];   // modexp_top.v(751)
    assign n7669 = rst ? encrypted_data_buf[1994] : encrypted_data_buf_next[1994];   // modexp_top.v(751)
    assign n7670 = rst ? encrypted_data_buf[1993] : encrypted_data_buf_next[1993];   // modexp_top.v(751)
    assign n7671 = rst ? encrypted_data_buf[1992] : encrypted_data_buf_next[1992];   // modexp_top.v(751)
    assign n7672 = rst ? encrypted_data_buf[1991] : encrypted_data_buf_next[1991];   // modexp_top.v(751)
    assign n7673 = rst ? encrypted_data_buf[1990] : encrypted_data_buf_next[1990];   // modexp_top.v(751)
    assign n7674 = rst ? encrypted_data_buf[1989] : encrypted_data_buf_next[1989];   // modexp_top.v(751)
    assign n7675 = rst ? encrypted_data_buf[1988] : encrypted_data_buf_next[1988];   // modexp_top.v(751)
    assign n7676 = rst ? encrypted_data_buf[1987] : encrypted_data_buf_next[1987];   // modexp_top.v(751)
    assign n7677 = rst ? encrypted_data_buf[1986] : encrypted_data_buf_next[1986];   // modexp_top.v(751)
    assign n7678 = rst ? encrypted_data_buf[1985] : encrypted_data_buf_next[1985];   // modexp_top.v(751)
    assign n7679 = rst ? encrypted_data_buf[1984] : encrypted_data_buf_next[1984];   // modexp_top.v(751)
    assign n7680 = rst ? encrypted_data_buf[1983] : encrypted_data_buf_next[1983];   // modexp_top.v(751)
    assign n7681 = rst ? encrypted_data_buf[1982] : encrypted_data_buf_next[1982];   // modexp_top.v(751)
    assign n7682 = rst ? encrypted_data_buf[1981] : encrypted_data_buf_next[1981];   // modexp_top.v(751)
    assign n7683 = rst ? encrypted_data_buf[1980] : encrypted_data_buf_next[1980];   // modexp_top.v(751)
    assign n7684 = rst ? encrypted_data_buf[1979] : encrypted_data_buf_next[1979];   // modexp_top.v(751)
    assign n7685 = rst ? encrypted_data_buf[1978] : encrypted_data_buf_next[1978];   // modexp_top.v(751)
    assign n7686 = rst ? encrypted_data_buf[1977] : encrypted_data_buf_next[1977];   // modexp_top.v(751)
    assign n7687 = rst ? encrypted_data_buf[1976] : encrypted_data_buf_next[1976];   // modexp_top.v(751)
    assign n7688 = rst ? encrypted_data_buf[1975] : encrypted_data_buf_next[1975];   // modexp_top.v(751)
    assign n7689 = rst ? encrypted_data_buf[1974] : encrypted_data_buf_next[1974];   // modexp_top.v(751)
    assign n7690 = rst ? encrypted_data_buf[1973] : encrypted_data_buf_next[1973];   // modexp_top.v(751)
    assign n7691 = rst ? encrypted_data_buf[1972] : encrypted_data_buf_next[1972];   // modexp_top.v(751)
    assign n7692 = rst ? encrypted_data_buf[1971] : encrypted_data_buf_next[1971];   // modexp_top.v(751)
    assign n7693 = rst ? encrypted_data_buf[1970] : encrypted_data_buf_next[1970];   // modexp_top.v(751)
    assign n7694 = rst ? encrypted_data_buf[1969] : encrypted_data_buf_next[1969];   // modexp_top.v(751)
    assign n7695 = rst ? encrypted_data_buf[1968] : encrypted_data_buf_next[1968];   // modexp_top.v(751)
    assign n7696 = rst ? encrypted_data_buf[1967] : encrypted_data_buf_next[1967];   // modexp_top.v(751)
    assign n7697 = rst ? encrypted_data_buf[1966] : encrypted_data_buf_next[1966];   // modexp_top.v(751)
    assign n7698 = rst ? encrypted_data_buf[1965] : encrypted_data_buf_next[1965];   // modexp_top.v(751)
    assign n7699 = rst ? encrypted_data_buf[1964] : encrypted_data_buf_next[1964];   // modexp_top.v(751)
    assign n7700 = rst ? encrypted_data_buf[1963] : encrypted_data_buf_next[1963];   // modexp_top.v(751)
    assign n7701 = rst ? encrypted_data_buf[1962] : encrypted_data_buf_next[1962];   // modexp_top.v(751)
    assign n7702 = rst ? encrypted_data_buf[1961] : encrypted_data_buf_next[1961];   // modexp_top.v(751)
    assign n7703 = rst ? encrypted_data_buf[1960] : encrypted_data_buf_next[1960];   // modexp_top.v(751)
    assign n7704 = rst ? encrypted_data_buf[1959] : encrypted_data_buf_next[1959];   // modexp_top.v(751)
    assign n7705 = rst ? encrypted_data_buf[1958] : encrypted_data_buf_next[1958];   // modexp_top.v(751)
    assign n7706 = rst ? encrypted_data_buf[1957] : encrypted_data_buf_next[1957];   // modexp_top.v(751)
    assign n7707 = rst ? encrypted_data_buf[1956] : encrypted_data_buf_next[1956];   // modexp_top.v(751)
    assign n7708 = rst ? encrypted_data_buf[1955] : encrypted_data_buf_next[1955];   // modexp_top.v(751)
    assign n7709 = rst ? encrypted_data_buf[1954] : encrypted_data_buf_next[1954];   // modexp_top.v(751)
    assign n7710 = rst ? encrypted_data_buf[1953] : encrypted_data_buf_next[1953];   // modexp_top.v(751)
    assign n7711 = rst ? encrypted_data_buf[1952] : encrypted_data_buf_next[1952];   // modexp_top.v(751)
    assign n7712 = rst ? encrypted_data_buf[1951] : encrypted_data_buf_next[1951];   // modexp_top.v(751)
    assign n7713 = rst ? encrypted_data_buf[1950] : encrypted_data_buf_next[1950];   // modexp_top.v(751)
    assign n7714 = rst ? encrypted_data_buf[1949] : encrypted_data_buf_next[1949];   // modexp_top.v(751)
    assign n7715 = rst ? encrypted_data_buf[1948] : encrypted_data_buf_next[1948];   // modexp_top.v(751)
    assign n7716 = rst ? encrypted_data_buf[1947] : encrypted_data_buf_next[1947];   // modexp_top.v(751)
    assign n7717 = rst ? encrypted_data_buf[1946] : encrypted_data_buf_next[1946];   // modexp_top.v(751)
    assign n7718 = rst ? encrypted_data_buf[1945] : encrypted_data_buf_next[1945];   // modexp_top.v(751)
    assign n7719 = rst ? encrypted_data_buf[1944] : encrypted_data_buf_next[1944];   // modexp_top.v(751)
    assign n7720 = rst ? encrypted_data_buf[1943] : encrypted_data_buf_next[1943];   // modexp_top.v(751)
    assign n7721 = rst ? encrypted_data_buf[1942] : encrypted_data_buf_next[1942];   // modexp_top.v(751)
    assign n7722 = rst ? encrypted_data_buf[1941] : encrypted_data_buf_next[1941];   // modexp_top.v(751)
    assign n7723 = rst ? encrypted_data_buf[1940] : encrypted_data_buf_next[1940];   // modexp_top.v(751)
    assign n7724 = rst ? encrypted_data_buf[1939] : encrypted_data_buf_next[1939];   // modexp_top.v(751)
    assign n7725 = rst ? encrypted_data_buf[1938] : encrypted_data_buf_next[1938];   // modexp_top.v(751)
    assign n7726 = rst ? encrypted_data_buf[1937] : encrypted_data_buf_next[1937];   // modexp_top.v(751)
    assign n7727 = rst ? encrypted_data_buf[1936] : encrypted_data_buf_next[1936];   // modexp_top.v(751)
    assign n7728 = rst ? encrypted_data_buf[1935] : encrypted_data_buf_next[1935];   // modexp_top.v(751)
    assign n7729 = rst ? encrypted_data_buf[1934] : encrypted_data_buf_next[1934];   // modexp_top.v(751)
    assign n7730 = rst ? encrypted_data_buf[1933] : encrypted_data_buf_next[1933];   // modexp_top.v(751)
    assign n7731 = rst ? encrypted_data_buf[1932] : encrypted_data_buf_next[1932];   // modexp_top.v(751)
    assign n7732 = rst ? encrypted_data_buf[1931] : encrypted_data_buf_next[1931];   // modexp_top.v(751)
    assign n7733 = rst ? encrypted_data_buf[1930] : encrypted_data_buf_next[1930];   // modexp_top.v(751)
    assign n7734 = rst ? encrypted_data_buf[1929] : encrypted_data_buf_next[1929];   // modexp_top.v(751)
    assign n7735 = rst ? encrypted_data_buf[1928] : encrypted_data_buf_next[1928];   // modexp_top.v(751)
    assign n7736 = rst ? encrypted_data_buf[1927] : encrypted_data_buf_next[1927];   // modexp_top.v(751)
    assign n7737 = rst ? encrypted_data_buf[1926] : encrypted_data_buf_next[1926];   // modexp_top.v(751)
    assign n7738 = rst ? encrypted_data_buf[1925] : encrypted_data_buf_next[1925];   // modexp_top.v(751)
    assign n7739 = rst ? encrypted_data_buf[1924] : encrypted_data_buf_next[1924];   // modexp_top.v(751)
    assign n7740 = rst ? encrypted_data_buf[1923] : encrypted_data_buf_next[1923];   // modexp_top.v(751)
    assign n7741 = rst ? encrypted_data_buf[1922] : encrypted_data_buf_next[1922];   // modexp_top.v(751)
    assign n7742 = rst ? encrypted_data_buf[1921] : encrypted_data_buf_next[1921];   // modexp_top.v(751)
    assign n7743 = rst ? encrypted_data_buf[1920] : encrypted_data_buf_next[1920];   // modexp_top.v(751)
    assign n7744 = rst ? encrypted_data_buf[1919] : encrypted_data_buf_next[1919];   // modexp_top.v(751)
    assign n7745 = rst ? encrypted_data_buf[1918] : encrypted_data_buf_next[1918];   // modexp_top.v(751)
    assign n7746 = rst ? encrypted_data_buf[1917] : encrypted_data_buf_next[1917];   // modexp_top.v(751)
    assign n7747 = rst ? encrypted_data_buf[1916] : encrypted_data_buf_next[1916];   // modexp_top.v(751)
    assign n7748 = rst ? encrypted_data_buf[1915] : encrypted_data_buf_next[1915];   // modexp_top.v(751)
    assign n7749 = rst ? encrypted_data_buf[1914] : encrypted_data_buf_next[1914];   // modexp_top.v(751)
    assign n7750 = rst ? encrypted_data_buf[1913] : encrypted_data_buf_next[1913];   // modexp_top.v(751)
    assign n7751 = rst ? encrypted_data_buf[1912] : encrypted_data_buf_next[1912];   // modexp_top.v(751)
    assign n7752 = rst ? encrypted_data_buf[1911] : encrypted_data_buf_next[1911];   // modexp_top.v(751)
    assign n7753 = rst ? encrypted_data_buf[1910] : encrypted_data_buf_next[1910];   // modexp_top.v(751)
    assign n7754 = rst ? encrypted_data_buf[1909] : encrypted_data_buf_next[1909];   // modexp_top.v(751)
    assign n7755 = rst ? encrypted_data_buf[1908] : encrypted_data_buf_next[1908];   // modexp_top.v(751)
    assign n7756 = rst ? encrypted_data_buf[1907] : encrypted_data_buf_next[1907];   // modexp_top.v(751)
    assign n7757 = rst ? encrypted_data_buf[1906] : encrypted_data_buf_next[1906];   // modexp_top.v(751)
    assign n7758 = rst ? encrypted_data_buf[1905] : encrypted_data_buf_next[1905];   // modexp_top.v(751)
    assign n7759 = rst ? encrypted_data_buf[1904] : encrypted_data_buf_next[1904];   // modexp_top.v(751)
    assign n7760 = rst ? encrypted_data_buf[1903] : encrypted_data_buf_next[1903];   // modexp_top.v(751)
    assign n7761 = rst ? encrypted_data_buf[1902] : encrypted_data_buf_next[1902];   // modexp_top.v(751)
    assign n7762 = rst ? encrypted_data_buf[1901] : encrypted_data_buf_next[1901];   // modexp_top.v(751)
    assign n7763 = rst ? encrypted_data_buf[1900] : encrypted_data_buf_next[1900];   // modexp_top.v(751)
    assign n7764 = rst ? encrypted_data_buf[1899] : encrypted_data_buf_next[1899];   // modexp_top.v(751)
    assign n7765 = rst ? encrypted_data_buf[1898] : encrypted_data_buf_next[1898];   // modexp_top.v(751)
    assign n7766 = rst ? encrypted_data_buf[1897] : encrypted_data_buf_next[1897];   // modexp_top.v(751)
    assign n7767 = rst ? encrypted_data_buf[1896] : encrypted_data_buf_next[1896];   // modexp_top.v(751)
    assign n7768 = rst ? encrypted_data_buf[1895] : encrypted_data_buf_next[1895];   // modexp_top.v(751)
    assign n7769 = rst ? encrypted_data_buf[1894] : encrypted_data_buf_next[1894];   // modexp_top.v(751)
    assign n7770 = rst ? encrypted_data_buf[1893] : encrypted_data_buf_next[1893];   // modexp_top.v(751)
    assign n7771 = rst ? encrypted_data_buf[1892] : encrypted_data_buf_next[1892];   // modexp_top.v(751)
    assign n7772 = rst ? encrypted_data_buf[1891] : encrypted_data_buf_next[1891];   // modexp_top.v(751)
    assign n7773 = rst ? encrypted_data_buf[1890] : encrypted_data_buf_next[1890];   // modexp_top.v(751)
    assign n7774 = rst ? encrypted_data_buf[1889] : encrypted_data_buf_next[1889];   // modexp_top.v(751)
    assign n7775 = rst ? encrypted_data_buf[1888] : encrypted_data_buf_next[1888];   // modexp_top.v(751)
    assign n7776 = rst ? encrypted_data_buf[1887] : encrypted_data_buf_next[1887];   // modexp_top.v(751)
    assign n7777 = rst ? encrypted_data_buf[1886] : encrypted_data_buf_next[1886];   // modexp_top.v(751)
    assign n7778 = rst ? encrypted_data_buf[1885] : encrypted_data_buf_next[1885];   // modexp_top.v(751)
    assign n7779 = rst ? encrypted_data_buf[1884] : encrypted_data_buf_next[1884];   // modexp_top.v(751)
    assign n7780 = rst ? encrypted_data_buf[1883] : encrypted_data_buf_next[1883];   // modexp_top.v(751)
    assign n7781 = rst ? encrypted_data_buf[1882] : encrypted_data_buf_next[1882];   // modexp_top.v(751)
    assign n7782 = rst ? encrypted_data_buf[1881] : encrypted_data_buf_next[1881];   // modexp_top.v(751)
    assign n7783 = rst ? encrypted_data_buf[1880] : encrypted_data_buf_next[1880];   // modexp_top.v(751)
    assign n7784 = rst ? encrypted_data_buf[1879] : encrypted_data_buf_next[1879];   // modexp_top.v(751)
    assign n7785 = rst ? encrypted_data_buf[1878] : encrypted_data_buf_next[1878];   // modexp_top.v(751)
    assign n7786 = rst ? encrypted_data_buf[1877] : encrypted_data_buf_next[1877];   // modexp_top.v(751)
    assign n7787 = rst ? encrypted_data_buf[1876] : encrypted_data_buf_next[1876];   // modexp_top.v(751)
    assign n7788 = rst ? encrypted_data_buf[1875] : encrypted_data_buf_next[1875];   // modexp_top.v(751)
    assign n7789 = rst ? encrypted_data_buf[1874] : encrypted_data_buf_next[1874];   // modexp_top.v(751)
    assign n7790 = rst ? encrypted_data_buf[1873] : encrypted_data_buf_next[1873];   // modexp_top.v(751)
    assign n7791 = rst ? encrypted_data_buf[1872] : encrypted_data_buf_next[1872];   // modexp_top.v(751)
    assign n7792 = rst ? encrypted_data_buf[1871] : encrypted_data_buf_next[1871];   // modexp_top.v(751)
    assign n7793 = rst ? encrypted_data_buf[1870] : encrypted_data_buf_next[1870];   // modexp_top.v(751)
    assign n7794 = rst ? encrypted_data_buf[1869] : encrypted_data_buf_next[1869];   // modexp_top.v(751)
    assign n7795 = rst ? encrypted_data_buf[1868] : encrypted_data_buf_next[1868];   // modexp_top.v(751)
    assign n7796 = rst ? encrypted_data_buf[1867] : encrypted_data_buf_next[1867];   // modexp_top.v(751)
    assign n7797 = rst ? encrypted_data_buf[1866] : encrypted_data_buf_next[1866];   // modexp_top.v(751)
    assign n7798 = rst ? encrypted_data_buf[1865] : encrypted_data_buf_next[1865];   // modexp_top.v(751)
    assign n7799 = rst ? encrypted_data_buf[1864] : encrypted_data_buf_next[1864];   // modexp_top.v(751)
    assign n7800 = rst ? encrypted_data_buf[1863] : encrypted_data_buf_next[1863];   // modexp_top.v(751)
    assign n7801 = rst ? encrypted_data_buf[1862] : encrypted_data_buf_next[1862];   // modexp_top.v(751)
    assign n7802 = rst ? encrypted_data_buf[1861] : encrypted_data_buf_next[1861];   // modexp_top.v(751)
    assign n7803 = rst ? encrypted_data_buf[1860] : encrypted_data_buf_next[1860];   // modexp_top.v(751)
    assign n7804 = rst ? encrypted_data_buf[1859] : encrypted_data_buf_next[1859];   // modexp_top.v(751)
    assign n7805 = rst ? encrypted_data_buf[1858] : encrypted_data_buf_next[1858];   // modexp_top.v(751)
    assign n7806 = rst ? encrypted_data_buf[1857] : encrypted_data_buf_next[1857];   // modexp_top.v(751)
    assign n7807 = rst ? encrypted_data_buf[1856] : encrypted_data_buf_next[1856];   // modexp_top.v(751)
    assign n7808 = rst ? encrypted_data_buf[1855] : encrypted_data_buf_next[1855];   // modexp_top.v(751)
    assign n7809 = rst ? encrypted_data_buf[1854] : encrypted_data_buf_next[1854];   // modexp_top.v(751)
    assign n7810 = rst ? encrypted_data_buf[1853] : encrypted_data_buf_next[1853];   // modexp_top.v(751)
    assign n7811 = rst ? encrypted_data_buf[1852] : encrypted_data_buf_next[1852];   // modexp_top.v(751)
    assign n7812 = rst ? encrypted_data_buf[1851] : encrypted_data_buf_next[1851];   // modexp_top.v(751)
    assign n7813 = rst ? encrypted_data_buf[1850] : encrypted_data_buf_next[1850];   // modexp_top.v(751)
    assign n7814 = rst ? encrypted_data_buf[1849] : encrypted_data_buf_next[1849];   // modexp_top.v(751)
    assign n7815 = rst ? encrypted_data_buf[1848] : encrypted_data_buf_next[1848];   // modexp_top.v(751)
    assign n7816 = rst ? encrypted_data_buf[1847] : encrypted_data_buf_next[1847];   // modexp_top.v(751)
    assign n7817 = rst ? encrypted_data_buf[1846] : encrypted_data_buf_next[1846];   // modexp_top.v(751)
    assign n7818 = rst ? encrypted_data_buf[1845] : encrypted_data_buf_next[1845];   // modexp_top.v(751)
    assign n7819 = rst ? encrypted_data_buf[1844] : encrypted_data_buf_next[1844];   // modexp_top.v(751)
    assign n7820 = rst ? encrypted_data_buf[1843] : encrypted_data_buf_next[1843];   // modexp_top.v(751)
    assign n7821 = rst ? encrypted_data_buf[1842] : encrypted_data_buf_next[1842];   // modexp_top.v(751)
    assign n7822 = rst ? encrypted_data_buf[1841] : encrypted_data_buf_next[1841];   // modexp_top.v(751)
    assign n7823 = rst ? encrypted_data_buf[1840] : encrypted_data_buf_next[1840];   // modexp_top.v(751)
    assign n7824 = rst ? encrypted_data_buf[1839] : encrypted_data_buf_next[1839];   // modexp_top.v(751)
    assign n7825 = rst ? encrypted_data_buf[1838] : encrypted_data_buf_next[1838];   // modexp_top.v(751)
    assign n7826 = rst ? encrypted_data_buf[1837] : encrypted_data_buf_next[1837];   // modexp_top.v(751)
    assign n7827 = rst ? encrypted_data_buf[1836] : encrypted_data_buf_next[1836];   // modexp_top.v(751)
    assign n7828 = rst ? encrypted_data_buf[1835] : encrypted_data_buf_next[1835];   // modexp_top.v(751)
    assign n7829 = rst ? encrypted_data_buf[1834] : encrypted_data_buf_next[1834];   // modexp_top.v(751)
    assign n7830 = rst ? encrypted_data_buf[1833] : encrypted_data_buf_next[1833];   // modexp_top.v(751)
    assign n7831 = rst ? encrypted_data_buf[1832] : encrypted_data_buf_next[1832];   // modexp_top.v(751)
    assign n7832 = rst ? encrypted_data_buf[1831] : encrypted_data_buf_next[1831];   // modexp_top.v(751)
    assign n7833 = rst ? encrypted_data_buf[1830] : encrypted_data_buf_next[1830];   // modexp_top.v(751)
    assign n7834 = rst ? encrypted_data_buf[1829] : encrypted_data_buf_next[1829];   // modexp_top.v(751)
    assign n7835 = rst ? encrypted_data_buf[1828] : encrypted_data_buf_next[1828];   // modexp_top.v(751)
    assign n7836 = rst ? encrypted_data_buf[1827] : encrypted_data_buf_next[1827];   // modexp_top.v(751)
    assign n7837 = rst ? encrypted_data_buf[1826] : encrypted_data_buf_next[1826];   // modexp_top.v(751)
    assign n7838 = rst ? encrypted_data_buf[1825] : encrypted_data_buf_next[1825];   // modexp_top.v(751)
    assign n7839 = rst ? encrypted_data_buf[1824] : encrypted_data_buf_next[1824];   // modexp_top.v(751)
    assign n7840 = rst ? encrypted_data_buf[1823] : encrypted_data_buf_next[1823];   // modexp_top.v(751)
    assign n7841 = rst ? encrypted_data_buf[1822] : encrypted_data_buf_next[1822];   // modexp_top.v(751)
    assign n7842 = rst ? encrypted_data_buf[1821] : encrypted_data_buf_next[1821];   // modexp_top.v(751)
    assign n7843 = rst ? encrypted_data_buf[1820] : encrypted_data_buf_next[1820];   // modexp_top.v(751)
    assign n7844 = rst ? encrypted_data_buf[1819] : encrypted_data_buf_next[1819];   // modexp_top.v(751)
    assign n7845 = rst ? encrypted_data_buf[1818] : encrypted_data_buf_next[1818];   // modexp_top.v(751)
    assign n7846 = rst ? encrypted_data_buf[1817] : encrypted_data_buf_next[1817];   // modexp_top.v(751)
    assign n7847 = rst ? encrypted_data_buf[1816] : encrypted_data_buf_next[1816];   // modexp_top.v(751)
    assign n7848 = rst ? encrypted_data_buf[1815] : encrypted_data_buf_next[1815];   // modexp_top.v(751)
    assign n7849 = rst ? encrypted_data_buf[1814] : encrypted_data_buf_next[1814];   // modexp_top.v(751)
    assign n7850 = rst ? encrypted_data_buf[1813] : encrypted_data_buf_next[1813];   // modexp_top.v(751)
    assign n7851 = rst ? encrypted_data_buf[1812] : encrypted_data_buf_next[1812];   // modexp_top.v(751)
    assign n7852 = rst ? encrypted_data_buf[1811] : encrypted_data_buf_next[1811];   // modexp_top.v(751)
    assign n7853 = rst ? encrypted_data_buf[1810] : encrypted_data_buf_next[1810];   // modexp_top.v(751)
    assign n7854 = rst ? encrypted_data_buf[1809] : encrypted_data_buf_next[1809];   // modexp_top.v(751)
    assign n7855 = rst ? encrypted_data_buf[1808] : encrypted_data_buf_next[1808];   // modexp_top.v(751)
    assign n7856 = rst ? encrypted_data_buf[1807] : encrypted_data_buf_next[1807];   // modexp_top.v(751)
    assign n7857 = rst ? encrypted_data_buf[1806] : encrypted_data_buf_next[1806];   // modexp_top.v(751)
    assign n7858 = rst ? encrypted_data_buf[1805] : encrypted_data_buf_next[1805];   // modexp_top.v(751)
    assign n7859 = rst ? encrypted_data_buf[1804] : encrypted_data_buf_next[1804];   // modexp_top.v(751)
    assign n7860 = rst ? encrypted_data_buf[1803] : encrypted_data_buf_next[1803];   // modexp_top.v(751)
    assign n7861 = rst ? encrypted_data_buf[1802] : encrypted_data_buf_next[1802];   // modexp_top.v(751)
    assign n7862 = rst ? encrypted_data_buf[1801] : encrypted_data_buf_next[1801];   // modexp_top.v(751)
    assign n7863 = rst ? encrypted_data_buf[1800] : encrypted_data_buf_next[1800];   // modexp_top.v(751)
    assign n7864 = rst ? encrypted_data_buf[1799] : encrypted_data_buf_next[1799];   // modexp_top.v(751)
    assign n7865 = rst ? encrypted_data_buf[1798] : encrypted_data_buf_next[1798];   // modexp_top.v(751)
    assign n7866 = rst ? encrypted_data_buf[1797] : encrypted_data_buf_next[1797];   // modexp_top.v(751)
    assign n7867 = rst ? encrypted_data_buf[1796] : encrypted_data_buf_next[1796];   // modexp_top.v(751)
    assign n7868 = rst ? encrypted_data_buf[1795] : encrypted_data_buf_next[1795];   // modexp_top.v(751)
    assign n7869 = rst ? encrypted_data_buf[1794] : encrypted_data_buf_next[1794];   // modexp_top.v(751)
    assign n7870 = rst ? encrypted_data_buf[1793] : encrypted_data_buf_next[1793];   // modexp_top.v(751)
    assign n7871 = rst ? encrypted_data_buf[1792] : encrypted_data_buf_next[1792];   // modexp_top.v(751)
    assign n7872 = rst ? encrypted_data_buf[1791] : encrypted_data_buf_next[1791];   // modexp_top.v(751)
    assign n7873 = rst ? encrypted_data_buf[1790] : encrypted_data_buf_next[1790];   // modexp_top.v(751)
    assign n7874 = rst ? encrypted_data_buf[1789] : encrypted_data_buf_next[1789];   // modexp_top.v(751)
    assign n7875 = rst ? encrypted_data_buf[1788] : encrypted_data_buf_next[1788];   // modexp_top.v(751)
    assign n7876 = rst ? encrypted_data_buf[1787] : encrypted_data_buf_next[1787];   // modexp_top.v(751)
    assign n7877 = rst ? encrypted_data_buf[1786] : encrypted_data_buf_next[1786];   // modexp_top.v(751)
    assign n7878 = rst ? encrypted_data_buf[1785] : encrypted_data_buf_next[1785];   // modexp_top.v(751)
    assign n7879 = rst ? encrypted_data_buf[1784] : encrypted_data_buf_next[1784];   // modexp_top.v(751)
    assign n7880 = rst ? encrypted_data_buf[1783] : encrypted_data_buf_next[1783];   // modexp_top.v(751)
    assign n7881 = rst ? encrypted_data_buf[1782] : encrypted_data_buf_next[1782];   // modexp_top.v(751)
    assign n7882 = rst ? encrypted_data_buf[1781] : encrypted_data_buf_next[1781];   // modexp_top.v(751)
    assign n7883 = rst ? encrypted_data_buf[1780] : encrypted_data_buf_next[1780];   // modexp_top.v(751)
    assign n7884 = rst ? encrypted_data_buf[1779] : encrypted_data_buf_next[1779];   // modexp_top.v(751)
    assign n7885 = rst ? encrypted_data_buf[1778] : encrypted_data_buf_next[1778];   // modexp_top.v(751)
    assign n7886 = rst ? encrypted_data_buf[1777] : encrypted_data_buf_next[1777];   // modexp_top.v(751)
    assign n7887 = rst ? encrypted_data_buf[1776] : encrypted_data_buf_next[1776];   // modexp_top.v(751)
    assign n7888 = rst ? encrypted_data_buf[1775] : encrypted_data_buf_next[1775];   // modexp_top.v(751)
    assign n7889 = rst ? encrypted_data_buf[1774] : encrypted_data_buf_next[1774];   // modexp_top.v(751)
    assign n7890 = rst ? encrypted_data_buf[1773] : encrypted_data_buf_next[1773];   // modexp_top.v(751)
    assign n7891 = rst ? encrypted_data_buf[1772] : encrypted_data_buf_next[1772];   // modexp_top.v(751)
    assign n7892 = rst ? encrypted_data_buf[1771] : encrypted_data_buf_next[1771];   // modexp_top.v(751)
    assign n7893 = rst ? encrypted_data_buf[1770] : encrypted_data_buf_next[1770];   // modexp_top.v(751)
    assign n7894 = rst ? encrypted_data_buf[1769] : encrypted_data_buf_next[1769];   // modexp_top.v(751)
    assign n7895 = rst ? encrypted_data_buf[1768] : encrypted_data_buf_next[1768];   // modexp_top.v(751)
    assign n7896 = rst ? encrypted_data_buf[1767] : encrypted_data_buf_next[1767];   // modexp_top.v(751)
    assign n7897 = rst ? encrypted_data_buf[1766] : encrypted_data_buf_next[1766];   // modexp_top.v(751)
    assign n7898 = rst ? encrypted_data_buf[1765] : encrypted_data_buf_next[1765];   // modexp_top.v(751)
    assign n7899 = rst ? encrypted_data_buf[1764] : encrypted_data_buf_next[1764];   // modexp_top.v(751)
    assign n7900 = rst ? encrypted_data_buf[1763] : encrypted_data_buf_next[1763];   // modexp_top.v(751)
    assign n7901 = rst ? encrypted_data_buf[1762] : encrypted_data_buf_next[1762];   // modexp_top.v(751)
    assign n7902 = rst ? encrypted_data_buf[1761] : encrypted_data_buf_next[1761];   // modexp_top.v(751)
    assign n7903 = rst ? encrypted_data_buf[1760] : encrypted_data_buf_next[1760];   // modexp_top.v(751)
    assign n7904 = rst ? encrypted_data_buf[1759] : encrypted_data_buf_next[1759];   // modexp_top.v(751)
    assign n7905 = rst ? encrypted_data_buf[1758] : encrypted_data_buf_next[1758];   // modexp_top.v(751)
    assign n7906 = rst ? encrypted_data_buf[1757] : encrypted_data_buf_next[1757];   // modexp_top.v(751)
    assign n7907 = rst ? encrypted_data_buf[1756] : encrypted_data_buf_next[1756];   // modexp_top.v(751)
    assign n7908 = rst ? encrypted_data_buf[1755] : encrypted_data_buf_next[1755];   // modexp_top.v(751)
    assign n7909 = rst ? encrypted_data_buf[1754] : encrypted_data_buf_next[1754];   // modexp_top.v(751)
    assign n7910 = rst ? encrypted_data_buf[1753] : encrypted_data_buf_next[1753];   // modexp_top.v(751)
    assign n7911 = rst ? encrypted_data_buf[1752] : encrypted_data_buf_next[1752];   // modexp_top.v(751)
    assign n7912 = rst ? encrypted_data_buf[1751] : encrypted_data_buf_next[1751];   // modexp_top.v(751)
    assign n7913 = rst ? encrypted_data_buf[1750] : encrypted_data_buf_next[1750];   // modexp_top.v(751)
    assign n7914 = rst ? encrypted_data_buf[1749] : encrypted_data_buf_next[1749];   // modexp_top.v(751)
    assign n7915 = rst ? encrypted_data_buf[1748] : encrypted_data_buf_next[1748];   // modexp_top.v(751)
    assign n7916 = rst ? encrypted_data_buf[1747] : encrypted_data_buf_next[1747];   // modexp_top.v(751)
    assign n7917 = rst ? encrypted_data_buf[1746] : encrypted_data_buf_next[1746];   // modexp_top.v(751)
    assign n7918 = rst ? encrypted_data_buf[1745] : encrypted_data_buf_next[1745];   // modexp_top.v(751)
    assign n7919 = rst ? encrypted_data_buf[1744] : encrypted_data_buf_next[1744];   // modexp_top.v(751)
    assign n7920 = rst ? encrypted_data_buf[1743] : encrypted_data_buf_next[1743];   // modexp_top.v(751)
    assign n7921 = rst ? encrypted_data_buf[1742] : encrypted_data_buf_next[1742];   // modexp_top.v(751)
    assign n7922 = rst ? encrypted_data_buf[1741] : encrypted_data_buf_next[1741];   // modexp_top.v(751)
    assign n7923 = rst ? encrypted_data_buf[1740] : encrypted_data_buf_next[1740];   // modexp_top.v(751)
    assign n7924 = rst ? encrypted_data_buf[1739] : encrypted_data_buf_next[1739];   // modexp_top.v(751)
    assign n7925 = rst ? encrypted_data_buf[1738] : encrypted_data_buf_next[1738];   // modexp_top.v(751)
    assign n7926 = rst ? encrypted_data_buf[1737] : encrypted_data_buf_next[1737];   // modexp_top.v(751)
    assign n7927 = rst ? encrypted_data_buf[1736] : encrypted_data_buf_next[1736];   // modexp_top.v(751)
    assign n7928 = rst ? encrypted_data_buf[1735] : encrypted_data_buf_next[1735];   // modexp_top.v(751)
    assign n7929 = rst ? encrypted_data_buf[1734] : encrypted_data_buf_next[1734];   // modexp_top.v(751)
    assign n7930 = rst ? encrypted_data_buf[1733] : encrypted_data_buf_next[1733];   // modexp_top.v(751)
    assign n7931 = rst ? encrypted_data_buf[1732] : encrypted_data_buf_next[1732];   // modexp_top.v(751)
    assign n7932 = rst ? encrypted_data_buf[1731] : encrypted_data_buf_next[1731];   // modexp_top.v(751)
    assign n7933 = rst ? encrypted_data_buf[1730] : encrypted_data_buf_next[1730];   // modexp_top.v(751)
    assign n7934 = rst ? encrypted_data_buf[1729] : encrypted_data_buf_next[1729];   // modexp_top.v(751)
    assign n7935 = rst ? encrypted_data_buf[1728] : encrypted_data_buf_next[1728];   // modexp_top.v(751)
    assign n7936 = rst ? encrypted_data_buf[1727] : encrypted_data_buf_next[1727];   // modexp_top.v(751)
    assign n7937 = rst ? encrypted_data_buf[1726] : encrypted_data_buf_next[1726];   // modexp_top.v(751)
    assign n7938 = rst ? encrypted_data_buf[1725] : encrypted_data_buf_next[1725];   // modexp_top.v(751)
    assign n7939 = rst ? encrypted_data_buf[1724] : encrypted_data_buf_next[1724];   // modexp_top.v(751)
    assign n7940 = rst ? encrypted_data_buf[1723] : encrypted_data_buf_next[1723];   // modexp_top.v(751)
    assign n7941 = rst ? encrypted_data_buf[1722] : encrypted_data_buf_next[1722];   // modexp_top.v(751)
    assign n7942 = rst ? encrypted_data_buf[1721] : encrypted_data_buf_next[1721];   // modexp_top.v(751)
    assign n7943 = rst ? encrypted_data_buf[1720] : encrypted_data_buf_next[1720];   // modexp_top.v(751)
    assign n7944 = rst ? encrypted_data_buf[1719] : encrypted_data_buf_next[1719];   // modexp_top.v(751)
    assign n7945 = rst ? encrypted_data_buf[1718] : encrypted_data_buf_next[1718];   // modexp_top.v(751)
    assign n7946 = rst ? encrypted_data_buf[1717] : encrypted_data_buf_next[1717];   // modexp_top.v(751)
    assign n7947 = rst ? encrypted_data_buf[1716] : encrypted_data_buf_next[1716];   // modexp_top.v(751)
    assign n7948 = rst ? encrypted_data_buf[1715] : encrypted_data_buf_next[1715];   // modexp_top.v(751)
    assign n7949 = rst ? encrypted_data_buf[1714] : encrypted_data_buf_next[1714];   // modexp_top.v(751)
    assign n7950 = rst ? encrypted_data_buf[1713] : encrypted_data_buf_next[1713];   // modexp_top.v(751)
    assign n7951 = rst ? encrypted_data_buf[1712] : encrypted_data_buf_next[1712];   // modexp_top.v(751)
    assign n7952 = rst ? encrypted_data_buf[1711] : encrypted_data_buf_next[1711];   // modexp_top.v(751)
    assign n7953 = rst ? encrypted_data_buf[1710] : encrypted_data_buf_next[1710];   // modexp_top.v(751)
    assign n7954 = rst ? encrypted_data_buf[1709] : encrypted_data_buf_next[1709];   // modexp_top.v(751)
    assign n7955 = rst ? encrypted_data_buf[1708] : encrypted_data_buf_next[1708];   // modexp_top.v(751)
    assign n7956 = rst ? encrypted_data_buf[1707] : encrypted_data_buf_next[1707];   // modexp_top.v(751)
    assign n7957 = rst ? encrypted_data_buf[1706] : encrypted_data_buf_next[1706];   // modexp_top.v(751)
    assign n7958 = rst ? encrypted_data_buf[1705] : encrypted_data_buf_next[1705];   // modexp_top.v(751)
    assign n7959 = rst ? encrypted_data_buf[1704] : encrypted_data_buf_next[1704];   // modexp_top.v(751)
    assign n7960 = rst ? encrypted_data_buf[1703] : encrypted_data_buf_next[1703];   // modexp_top.v(751)
    assign n7961 = rst ? encrypted_data_buf[1702] : encrypted_data_buf_next[1702];   // modexp_top.v(751)
    assign n7962 = rst ? encrypted_data_buf[1701] : encrypted_data_buf_next[1701];   // modexp_top.v(751)
    assign n7963 = rst ? encrypted_data_buf[1700] : encrypted_data_buf_next[1700];   // modexp_top.v(751)
    assign n7964 = rst ? encrypted_data_buf[1699] : encrypted_data_buf_next[1699];   // modexp_top.v(751)
    assign n7965 = rst ? encrypted_data_buf[1698] : encrypted_data_buf_next[1698];   // modexp_top.v(751)
    assign n7966 = rst ? encrypted_data_buf[1697] : encrypted_data_buf_next[1697];   // modexp_top.v(751)
    assign n7967 = rst ? encrypted_data_buf[1696] : encrypted_data_buf_next[1696];   // modexp_top.v(751)
    assign n7968 = rst ? encrypted_data_buf[1695] : encrypted_data_buf_next[1695];   // modexp_top.v(751)
    assign n7969 = rst ? encrypted_data_buf[1694] : encrypted_data_buf_next[1694];   // modexp_top.v(751)
    assign n7970 = rst ? encrypted_data_buf[1693] : encrypted_data_buf_next[1693];   // modexp_top.v(751)
    assign n7971 = rst ? encrypted_data_buf[1692] : encrypted_data_buf_next[1692];   // modexp_top.v(751)
    assign n7972 = rst ? encrypted_data_buf[1691] : encrypted_data_buf_next[1691];   // modexp_top.v(751)
    assign n7973 = rst ? encrypted_data_buf[1690] : encrypted_data_buf_next[1690];   // modexp_top.v(751)
    assign n7974 = rst ? encrypted_data_buf[1689] : encrypted_data_buf_next[1689];   // modexp_top.v(751)
    assign n7975 = rst ? encrypted_data_buf[1688] : encrypted_data_buf_next[1688];   // modexp_top.v(751)
    assign n7976 = rst ? encrypted_data_buf[1687] : encrypted_data_buf_next[1687];   // modexp_top.v(751)
    assign n7977 = rst ? encrypted_data_buf[1686] : encrypted_data_buf_next[1686];   // modexp_top.v(751)
    assign n7978 = rst ? encrypted_data_buf[1685] : encrypted_data_buf_next[1685];   // modexp_top.v(751)
    assign n7979 = rst ? encrypted_data_buf[1684] : encrypted_data_buf_next[1684];   // modexp_top.v(751)
    assign n7980 = rst ? encrypted_data_buf[1683] : encrypted_data_buf_next[1683];   // modexp_top.v(751)
    assign n7981 = rst ? encrypted_data_buf[1682] : encrypted_data_buf_next[1682];   // modexp_top.v(751)
    assign n7982 = rst ? encrypted_data_buf[1681] : encrypted_data_buf_next[1681];   // modexp_top.v(751)
    assign n7983 = rst ? encrypted_data_buf[1680] : encrypted_data_buf_next[1680];   // modexp_top.v(751)
    assign n7984 = rst ? encrypted_data_buf[1679] : encrypted_data_buf_next[1679];   // modexp_top.v(751)
    assign n7985 = rst ? encrypted_data_buf[1678] : encrypted_data_buf_next[1678];   // modexp_top.v(751)
    assign n7986 = rst ? encrypted_data_buf[1677] : encrypted_data_buf_next[1677];   // modexp_top.v(751)
    assign n7987 = rst ? encrypted_data_buf[1676] : encrypted_data_buf_next[1676];   // modexp_top.v(751)
    assign n7988 = rst ? encrypted_data_buf[1675] : encrypted_data_buf_next[1675];   // modexp_top.v(751)
    assign n7989 = rst ? encrypted_data_buf[1674] : encrypted_data_buf_next[1674];   // modexp_top.v(751)
    assign n7990 = rst ? encrypted_data_buf[1673] : encrypted_data_buf_next[1673];   // modexp_top.v(751)
    assign n7991 = rst ? encrypted_data_buf[1672] : encrypted_data_buf_next[1672];   // modexp_top.v(751)
    assign n7992 = rst ? encrypted_data_buf[1671] : encrypted_data_buf_next[1671];   // modexp_top.v(751)
    assign n7993 = rst ? encrypted_data_buf[1670] : encrypted_data_buf_next[1670];   // modexp_top.v(751)
    assign n7994 = rst ? encrypted_data_buf[1669] : encrypted_data_buf_next[1669];   // modexp_top.v(751)
    assign n7995 = rst ? encrypted_data_buf[1668] : encrypted_data_buf_next[1668];   // modexp_top.v(751)
    assign n7996 = rst ? encrypted_data_buf[1667] : encrypted_data_buf_next[1667];   // modexp_top.v(751)
    assign n7997 = rst ? encrypted_data_buf[1666] : encrypted_data_buf_next[1666];   // modexp_top.v(751)
    assign n7998 = rst ? encrypted_data_buf[1665] : encrypted_data_buf_next[1665];   // modexp_top.v(751)
    assign n7999 = rst ? encrypted_data_buf[1664] : encrypted_data_buf_next[1664];   // modexp_top.v(751)
    assign n8000 = rst ? encrypted_data_buf[1663] : encrypted_data_buf_next[1663];   // modexp_top.v(751)
    assign n8001 = rst ? encrypted_data_buf[1662] : encrypted_data_buf_next[1662];   // modexp_top.v(751)
    assign n8002 = rst ? encrypted_data_buf[1661] : encrypted_data_buf_next[1661];   // modexp_top.v(751)
    assign n8003 = rst ? encrypted_data_buf[1660] : encrypted_data_buf_next[1660];   // modexp_top.v(751)
    assign n8004 = rst ? encrypted_data_buf[1659] : encrypted_data_buf_next[1659];   // modexp_top.v(751)
    assign n8005 = rst ? encrypted_data_buf[1658] : encrypted_data_buf_next[1658];   // modexp_top.v(751)
    assign n8006 = rst ? encrypted_data_buf[1657] : encrypted_data_buf_next[1657];   // modexp_top.v(751)
    assign n8007 = rst ? encrypted_data_buf[1656] : encrypted_data_buf_next[1656];   // modexp_top.v(751)
    assign n8008 = rst ? encrypted_data_buf[1655] : encrypted_data_buf_next[1655];   // modexp_top.v(751)
    assign n8009 = rst ? encrypted_data_buf[1654] : encrypted_data_buf_next[1654];   // modexp_top.v(751)
    assign n8010 = rst ? encrypted_data_buf[1653] : encrypted_data_buf_next[1653];   // modexp_top.v(751)
    assign n8011 = rst ? encrypted_data_buf[1652] : encrypted_data_buf_next[1652];   // modexp_top.v(751)
    assign n8012 = rst ? encrypted_data_buf[1651] : encrypted_data_buf_next[1651];   // modexp_top.v(751)
    assign n8013 = rst ? encrypted_data_buf[1650] : encrypted_data_buf_next[1650];   // modexp_top.v(751)
    assign n8014 = rst ? encrypted_data_buf[1649] : encrypted_data_buf_next[1649];   // modexp_top.v(751)
    assign n8015 = rst ? encrypted_data_buf[1648] : encrypted_data_buf_next[1648];   // modexp_top.v(751)
    assign n8016 = rst ? encrypted_data_buf[1647] : encrypted_data_buf_next[1647];   // modexp_top.v(751)
    assign n8017 = rst ? encrypted_data_buf[1646] : encrypted_data_buf_next[1646];   // modexp_top.v(751)
    assign n8018 = rst ? encrypted_data_buf[1645] : encrypted_data_buf_next[1645];   // modexp_top.v(751)
    assign n8019 = rst ? encrypted_data_buf[1644] : encrypted_data_buf_next[1644];   // modexp_top.v(751)
    assign n8020 = rst ? encrypted_data_buf[1643] : encrypted_data_buf_next[1643];   // modexp_top.v(751)
    assign n8021 = rst ? encrypted_data_buf[1642] : encrypted_data_buf_next[1642];   // modexp_top.v(751)
    assign n8022 = rst ? encrypted_data_buf[1641] : encrypted_data_buf_next[1641];   // modexp_top.v(751)
    assign n8023 = rst ? encrypted_data_buf[1640] : encrypted_data_buf_next[1640];   // modexp_top.v(751)
    assign n8024 = rst ? encrypted_data_buf[1639] : encrypted_data_buf_next[1639];   // modexp_top.v(751)
    assign n8025 = rst ? encrypted_data_buf[1638] : encrypted_data_buf_next[1638];   // modexp_top.v(751)
    assign n8026 = rst ? encrypted_data_buf[1637] : encrypted_data_buf_next[1637];   // modexp_top.v(751)
    assign n8027 = rst ? encrypted_data_buf[1636] : encrypted_data_buf_next[1636];   // modexp_top.v(751)
    assign n8028 = rst ? encrypted_data_buf[1635] : encrypted_data_buf_next[1635];   // modexp_top.v(751)
    assign n8029 = rst ? encrypted_data_buf[1634] : encrypted_data_buf_next[1634];   // modexp_top.v(751)
    assign n8030 = rst ? encrypted_data_buf[1633] : encrypted_data_buf_next[1633];   // modexp_top.v(751)
    assign n8031 = rst ? encrypted_data_buf[1632] : encrypted_data_buf_next[1632];   // modexp_top.v(751)
    assign n8032 = rst ? encrypted_data_buf[1631] : encrypted_data_buf_next[1631];   // modexp_top.v(751)
    assign n8033 = rst ? encrypted_data_buf[1630] : encrypted_data_buf_next[1630];   // modexp_top.v(751)
    assign n8034 = rst ? encrypted_data_buf[1629] : encrypted_data_buf_next[1629];   // modexp_top.v(751)
    assign n8035 = rst ? encrypted_data_buf[1628] : encrypted_data_buf_next[1628];   // modexp_top.v(751)
    assign n8036 = rst ? encrypted_data_buf[1627] : encrypted_data_buf_next[1627];   // modexp_top.v(751)
    assign n8037 = rst ? encrypted_data_buf[1626] : encrypted_data_buf_next[1626];   // modexp_top.v(751)
    assign n8038 = rst ? encrypted_data_buf[1625] : encrypted_data_buf_next[1625];   // modexp_top.v(751)
    assign n8039 = rst ? encrypted_data_buf[1624] : encrypted_data_buf_next[1624];   // modexp_top.v(751)
    assign n8040 = rst ? encrypted_data_buf[1623] : encrypted_data_buf_next[1623];   // modexp_top.v(751)
    assign n8041 = rst ? encrypted_data_buf[1622] : encrypted_data_buf_next[1622];   // modexp_top.v(751)
    assign n8042 = rst ? encrypted_data_buf[1621] : encrypted_data_buf_next[1621];   // modexp_top.v(751)
    assign n8043 = rst ? encrypted_data_buf[1620] : encrypted_data_buf_next[1620];   // modexp_top.v(751)
    assign n8044 = rst ? encrypted_data_buf[1619] : encrypted_data_buf_next[1619];   // modexp_top.v(751)
    assign n8045 = rst ? encrypted_data_buf[1618] : encrypted_data_buf_next[1618];   // modexp_top.v(751)
    assign n8046 = rst ? encrypted_data_buf[1617] : encrypted_data_buf_next[1617];   // modexp_top.v(751)
    assign n8047 = rst ? encrypted_data_buf[1616] : encrypted_data_buf_next[1616];   // modexp_top.v(751)
    assign n8048 = rst ? encrypted_data_buf[1615] : encrypted_data_buf_next[1615];   // modexp_top.v(751)
    assign n8049 = rst ? encrypted_data_buf[1614] : encrypted_data_buf_next[1614];   // modexp_top.v(751)
    assign n8050 = rst ? encrypted_data_buf[1613] : encrypted_data_buf_next[1613];   // modexp_top.v(751)
    assign n8051 = rst ? encrypted_data_buf[1612] : encrypted_data_buf_next[1612];   // modexp_top.v(751)
    assign n8052 = rst ? encrypted_data_buf[1611] : encrypted_data_buf_next[1611];   // modexp_top.v(751)
    assign n8053 = rst ? encrypted_data_buf[1610] : encrypted_data_buf_next[1610];   // modexp_top.v(751)
    assign n8054 = rst ? encrypted_data_buf[1609] : encrypted_data_buf_next[1609];   // modexp_top.v(751)
    assign n8055 = rst ? encrypted_data_buf[1608] : encrypted_data_buf_next[1608];   // modexp_top.v(751)
    assign n8056 = rst ? encrypted_data_buf[1607] : encrypted_data_buf_next[1607];   // modexp_top.v(751)
    assign n8057 = rst ? encrypted_data_buf[1606] : encrypted_data_buf_next[1606];   // modexp_top.v(751)
    assign n8058 = rst ? encrypted_data_buf[1605] : encrypted_data_buf_next[1605];   // modexp_top.v(751)
    assign n8059 = rst ? encrypted_data_buf[1604] : encrypted_data_buf_next[1604];   // modexp_top.v(751)
    assign n8060 = rst ? encrypted_data_buf[1603] : encrypted_data_buf_next[1603];   // modexp_top.v(751)
    assign n8061 = rst ? encrypted_data_buf[1602] : encrypted_data_buf_next[1602];   // modexp_top.v(751)
    assign n8062 = rst ? encrypted_data_buf[1601] : encrypted_data_buf_next[1601];   // modexp_top.v(751)
    assign n8063 = rst ? encrypted_data_buf[1600] : encrypted_data_buf_next[1600];   // modexp_top.v(751)
    assign n8064 = rst ? encrypted_data_buf[1599] : encrypted_data_buf_next[1599];   // modexp_top.v(751)
    assign n8065 = rst ? encrypted_data_buf[1598] : encrypted_data_buf_next[1598];   // modexp_top.v(751)
    assign n8066 = rst ? encrypted_data_buf[1597] : encrypted_data_buf_next[1597];   // modexp_top.v(751)
    assign n8067 = rst ? encrypted_data_buf[1596] : encrypted_data_buf_next[1596];   // modexp_top.v(751)
    assign n8068 = rst ? encrypted_data_buf[1595] : encrypted_data_buf_next[1595];   // modexp_top.v(751)
    assign n8069 = rst ? encrypted_data_buf[1594] : encrypted_data_buf_next[1594];   // modexp_top.v(751)
    assign n8070 = rst ? encrypted_data_buf[1593] : encrypted_data_buf_next[1593];   // modexp_top.v(751)
    assign n8071 = rst ? encrypted_data_buf[1592] : encrypted_data_buf_next[1592];   // modexp_top.v(751)
    assign n8072 = rst ? encrypted_data_buf[1591] : encrypted_data_buf_next[1591];   // modexp_top.v(751)
    assign n8073 = rst ? encrypted_data_buf[1590] : encrypted_data_buf_next[1590];   // modexp_top.v(751)
    assign n8074 = rst ? encrypted_data_buf[1589] : encrypted_data_buf_next[1589];   // modexp_top.v(751)
    assign n8075 = rst ? encrypted_data_buf[1588] : encrypted_data_buf_next[1588];   // modexp_top.v(751)
    assign n8076 = rst ? encrypted_data_buf[1587] : encrypted_data_buf_next[1587];   // modexp_top.v(751)
    assign n8077 = rst ? encrypted_data_buf[1586] : encrypted_data_buf_next[1586];   // modexp_top.v(751)
    assign n8078 = rst ? encrypted_data_buf[1585] : encrypted_data_buf_next[1585];   // modexp_top.v(751)
    assign n8079 = rst ? encrypted_data_buf[1584] : encrypted_data_buf_next[1584];   // modexp_top.v(751)
    assign n8080 = rst ? encrypted_data_buf[1583] : encrypted_data_buf_next[1583];   // modexp_top.v(751)
    assign n8081 = rst ? encrypted_data_buf[1582] : encrypted_data_buf_next[1582];   // modexp_top.v(751)
    assign n8082 = rst ? encrypted_data_buf[1581] : encrypted_data_buf_next[1581];   // modexp_top.v(751)
    assign n8083 = rst ? encrypted_data_buf[1580] : encrypted_data_buf_next[1580];   // modexp_top.v(751)
    assign n8084 = rst ? encrypted_data_buf[1579] : encrypted_data_buf_next[1579];   // modexp_top.v(751)
    assign n8085 = rst ? encrypted_data_buf[1578] : encrypted_data_buf_next[1578];   // modexp_top.v(751)
    assign n8086 = rst ? encrypted_data_buf[1577] : encrypted_data_buf_next[1577];   // modexp_top.v(751)
    assign n8087 = rst ? encrypted_data_buf[1576] : encrypted_data_buf_next[1576];   // modexp_top.v(751)
    assign n8088 = rst ? encrypted_data_buf[1575] : encrypted_data_buf_next[1575];   // modexp_top.v(751)
    assign n8089 = rst ? encrypted_data_buf[1574] : encrypted_data_buf_next[1574];   // modexp_top.v(751)
    assign n8090 = rst ? encrypted_data_buf[1573] : encrypted_data_buf_next[1573];   // modexp_top.v(751)
    assign n8091 = rst ? encrypted_data_buf[1572] : encrypted_data_buf_next[1572];   // modexp_top.v(751)
    assign n8092 = rst ? encrypted_data_buf[1571] : encrypted_data_buf_next[1571];   // modexp_top.v(751)
    assign n8093 = rst ? encrypted_data_buf[1570] : encrypted_data_buf_next[1570];   // modexp_top.v(751)
    assign n8094 = rst ? encrypted_data_buf[1569] : encrypted_data_buf_next[1569];   // modexp_top.v(751)
    assign n8095 = rst ? encrypted_data_buf[1568] : encrypted_data_buf_next[1568];   // modexp_top.v(751)
    assign n8096 = rst ? encrypted_data_buf[1567] : encrypted_data_buf_next[1567];   // modexp_top.v(751)
    assign n8097 = rst ? encrypted_data_buf[1566] : encrypted_data_buf_next[1566];   // modexp_top.v(751)
    assign n8098 = rst ? encrypted_data_buf[1565] : encrypted_data_buf_next[1565];   // modexp_top.v(751)
    assign n8099 = rst ? encrypted_data_buf[1564] : encrypted_data_buf_next[1564];   // modexp_top.v(751)
    assign n8100 = rst ? encrypted_data_buf[1563] : encrypted_data_buf_next[1563];   // modexp_top.v(751)
    assign n8101 = rst ? encrypted_data_buf[1562] : encrypted_data_buf_next[1562];   // modexp_top.v(751)
    assign n8102 = rst ? encrypted_data_buf[1561] : encrypted_data_buf_next[1561];   // modexp_top.v(751)
    assign n8103 = rst ? encrypted_data_buf[1560] : encrypted_data_buf_next[1560];   // modexp_top.v(751)
    assign n8104 = rst ? encrypted_data_buf[1559] : encrypted_data_buf_next[1559];   // modexp_top.v(751)
    assign n8105 = rst ? encrypted_data_buf[1558] : encrypted_data_buf_next[1558];   // modexp_top.v(751)
    assign n8106 = rst ? encrypted_data_buf[1557] : encrypted_data_buf_next[1557];   // modexp_top.v(751)
    assign n8107 = rst ? encrypted_data_buf[1556] : encrypted_data_buf_next[1556];   // modexp_top.v(751)
    assign n8108 = rst ? encrypted_data_buf[1555] : encrypted_data_buf_next[1555];   // modexp_top.v(751)
    assign n8109 = rst ? encrypted_data_buf[1554] : encrypted_data_buf_next[1554];   // modexp_top.v(751)
    assign n8110 = rst ? encrypted_data_buf[1553] : encrypted_data_buf_next[1553];   // modexp_top.v(751)
    assign n8111 = rst ? encrypted_data_buf[1552] : encrypted_data_buf_next[1552];   // modexp_top.v(751)
    assign n8112 = rst ? encrypted_data_buf[1551] : encrypted_data_buf_next[1551];   // modexp_top.v(751)
    assign n8113 = rst ? encrypted_data_buf[1550] : encrypted_data_buf_next[1550];   // modexp_top.v(751)
    assign n8114 = rst ? encrypted_data_buf[1549] : encrypted_data_buf_next[1549];   // modexp_top.v(751)
    assign n8115 = rst ? encrypted_data_buf[1548] : encrypted_data_buf_next[1548];   // modexp_top.v(751)
    assign n8116 = rst ? encrypted_data_buf[1547] : encrypted_data_buf_next[1547];   // modexp_top.v(751)
    assign n8117 = rst ? encrypted_data_buf[1546] : encrypted_data_buf_next[1546];   // modexp_top.v(751)
    assign n8118 = rst ? encrypted_data_buf[1545] : encrypted_data_buf_next[1545];   // modexp_top.v(751)
    assign n8119 = rst ? encrypted_data_buf[1544] : encrypted_data_buf_next[1544];   // modexp_top.v(751)
    assign n8120 = rst ? encrypted_data_buf[1543] : encrypted_data_buf_next[1543];   // modexp_top.v(751)
    assign n8121 = rst ? encrypted_data_buf[1542] : encrypted_data_buf_next[1542];   // modexp_top.v(751)
    assign n8122 = rst ? encrypted_data_buf[1541] : encrypted_data_buf_next[1541];   // modexp_top.v(751)
    assign n8123 = rst ? encrypted_data_buf[1540] : encrypted_data_buf_next[1540];   // modexp_top.v(751)
    assign n8124 = rst ? encrypted_data_buf[1539] : encrypted_data_buf_next[1539];   // modexp_top.v(751)
    assign n8125 = rst ? encrypted_data_buf[1538] : encrypted_data_buf_next[1538];   // modexp_top.v(751)
    assign n8126 = rst ? encrypted_data_buf[1537] : encrypted_data_buf_next[1537];   // modexp_top.v(751)
    assign n8127 = rst ? encrypted_data_buf[1536] : encrypted_data_buf_next[1536];   // modexp_top.v(751)
    assign n8128 = rst ? encrypted_data_buf[1535] : encrypted_data_buf_next[1535];   // modexp_top.v(751)
    assign n8129 = rst ? encrypted_data_buf[1534] : encrypted_data_buf_next[1534];   // modexp_top.v(751)
    assign n8130 = rst ? encrypted_data_buf[1533] : encrypted_data_buf_next[1533];   // modexp_top.v(751)
    assign n8131 = rst ? encrypted_data_buf[1532] : encrypted_data_buf_next[1532];   // modexp_top.v(751)
    assign n8132 = rst ? encrypted_data_buf[1531] : encrypted_data_buf_next[1531];   // modexp_top.v(751)
    assign n8133 = rst ? encrypted_data_buf[1530] : encrypted_data_buf_next[1530];   // modexp_top.v(751)
    assign n8134 = rst ? encrypted_data_buf[1529] : encrypted_data_buf_next[1529];   // modexp_top.v(751)
    assign n8135 = rst ? encrypted_data_buf[1528] : encrypted_data_buf_next[1528];   // modexp_top.v(751)
    assign n8136 = rst ? encrypted_data_buf[1527] : encrypted_data_buf_next[1527];   // modexp_top.v(751)
    assign n8137 = rst ? encrypted_data_buf[1526] : encrypted_data_buf_next[1526];   // modexp_top.v(751)
    assign n8138 = rst ? encrypted_data_buf[1525] : encrypted_data_buf_next[1525];   // modexp_top.v(751)
    assign n8139 = rst ? encrypted_data_buf[1524] : encrypted_data_buf_next[1524];   // modexp_top.v(751)
    assign n8140 = rst ? encrypted_data_buf[1523] : encrypted_data_buf_next[1523];   // modexp_top.v(751)
    assign n8141 = rst ? encrypted_data_buf[1522] : encrypted_data_buf_next[1522];   // modexp_top.v(751)
    assign n8142 = rst ? encrypted_data_buf[1521] : encrypted_data_buf_next[1521];   // modexp_top.v(751)
    assign n8143 = rst ? encrypted_data_buf[1520] : encrypted_data_buf_next[1520];   // modexp_top.v(751)
    assign n8144 = rst ? encrypted_data_buf[1519] : encrypted_data_buf_next[1519];   // modexp_top.v(751)
    assign n8145 = rst ? encrypted_data_buf[1518] : encrypted_data_buf_next[1518];   // modexp_top.v(751)
    assign n8146 = rst ? encrypted_data_buf[1517] : encrypted_data_buf_next[1517];   // modexp_top.v(751)
    assign n8147 = rst ? encrypted_data_buf[1516] : encrypted_data_buf_next[1516];   // modexp_top.v(751)
    assign n8148 = rst ? encrypted_data_buf[1515] : encrypted_data_buf_next[1515];   // modexp_top.v(751)
    assign n8149 = rst ? encrypted_data_buf[1514] : encrypted_data_buf_next[1514];   // modexp_top.v(751)
    assign n8150 = rst ? encrypted_data_buf[1513] : encrypted_data_buf_next[1513];   // modexp_top.v(751)
    assign n8151 = rst ? encrypted_data_buf[1512] : encrypted_data_buf_next[1512];   // modexp_top.v(751)
    assign n8152 = rst ? encrypted_data_buf[1511] : encrypted_data_buf_next[1511];   // modexp_top.v(751)
    assign n8153 = rst ? encrypted_data_buf[1510] : encrypted_data_buf_next[1510];   // modexp_top.v(751)
    assign n8154 = rst ? encrypted_data_buf[1509] : encrypted_data_buf_next[1509];   // modexp_top.v(751)
    assign n8155 = rst ? encrypted_data_buf[1508] : encrypted_data_buf_next[1508];   // modexp_top.v(751)
    assign n8156 = rst ? encrypted_data_buf[1507] : encrypted_data_buf_next[1507];   // modexp_top.v(751)
    assign n8157 = rst ? encrypted_data_buf[1506] : encrypted_data_buf_next[1506];   // modexp_top.v(751)
    assign n8158 = rst ? encrypted_data_buf[1505] : encrypted_data_buf_next[1505];   // modexp_top.v(751)
    assign n8159 = rst ? encrypted_data_buf[1504] : encrypted_data_buf_next[1504];   // modexp_top.v(751)
    assign n8160 = rst ? encrypted_data_buf[1503] : encrypted_data_buf_next[1503];   // modexp_top.v(751)
    assign n8161 = rst ? encrypted_data_buf[1502] : encrypted_data_buf_next[1502];   // modexp_top.v(751)
    assign n8162 = rst ? encrypted_data_buf[1501] : encrypted_data_buf_next[1501];   // modexp_top.v(751)
    assign n8163 = rst ? encrypted_data_buf[1500] : encrypted_data_buf_next[1500];   // modexp_top.v(751)
    assign n8164 = rst ? encrypted_data_buf[1499] : encrypted_data_buf_next[1499];   // modexp_top.v(751)
    assign n8165 = rst ? encrypted_data_buf[1498] : encrypted_data_buf_next[1498];   // modexp_top.v(751)
    assign n8166 = rst ? encrypted_data_buf[1497] : encrypted_data_buf_next[1497];   // modexp_top.v(751)
    assign n8167 = rst ? encrypted_data_buf[1496] : encrypted_data_buf_next[1496];   // modexp_top.v(751)
    assign n8168 = rst ? encrypted_data_buf[1495] : encrypted_data_buf_next[1495];   // modexp_top.v(751)
    assign n8169 = rst ? encrypted_data_buf[1494] : encrypted_data_buf_next[1494];   // modexp_top.v(751)
    assign n8170 = rst ? encrypted_data_buf[1493] : encrypted_data_buf_next[1493];   // modexp_top.v(751)
    assign n8171 = rst ? encrypted_data_buf[1492] : encrypted_data_buf_next[1492];   // modexp_top.v(751)
    assign n8172 = rst ? encrypted_data_buf[1491] : encrypted_data_buf_next[1491];   // modexp_top.v(751)
    assign n8173 = rst ? encrypted_data_buf[1490] : encrypted_data_buf_next[1490];   // modexp_top.v(751)
    assign n8174 = rst ? encrypted_data_buf[1489] : encrypted_data_buf_next[1489];   // modexp_top.v(751)
    assign n8175 = rst ? encrypted_data_buf[1488] : encrypted_data_buf_next[1488];   // modexp_top.v(751)
    assign n8176 = rst ? encrypted_data_buf[1487] : encrypted_data_buf_next[1487];   // modexp_top.v(751)
    assign n8177 = rst ? encrypted_data_buf[1486] : encrypted_data_buf_next[1486];   // modexp_top.v(751)
    assign n8178 = rst ? encrypted_data_buf[1485] : encrypted_data_buf_next[1485];   // modexp_top.v(751)
    assign n8179 = rst ? encrypted_data_buf[1484] : encrypted_data_buf_next[1484];   // modexp_top.v(751)
    assign n8180 = rst ? encrypted_data_buf[1483] : encrypted_data_buf_next[1483];   // modexp_top.v(751)
    assign n8181 = rst ? encrypted_data_buf[1482] : encrypted_data_buf_next[1482];   // modexp_top.v(751)
    assign n8182 = rst ? encrypted_data_buf[1481] : encrypted_data_buf_next[1481];   // modexp_top.v(751)
    assign n8183 = rst ? encrypted_data_buf[1480] : encrypted_data_buf_next[1480];   // modexp_top.v(751)
    assign n8184 = rst ? encrypted_data_buf[1479] : encrypted_data_buf_next[1479];   // modexp_top.v(751)
    assign n8185 = rst ? encrypted_data_buf[1478] : encrypted_data_buf_next[1478];   // modexp_top.v(751)
    assign n8186 = rst ? encrypted_data_buf[1477] : encrypted_data_buf_next[1477];   // modexp_top.v(751)
    assign n8187 = rst ? encrypted_data_buf[1476] : encrypted_data_buf_next[1476];   // modexp_top.v(751)
    assign n8188 = rst ? encrypted_data_buf[1475] : encrypted_data_buf_next[1475];   // modexp_top.v(751)
    assign n8189 = rst ? encrypted_data_buf[1474] : encrypted_data_buf_next[1474];   // modexp_top.v(751)
    assign n8190 = rst ? encrypted_data_buf[1473] : encrypted_data_buf_next[1473];   // modexp_top.v(751)
    assign n8191 = rst ? encrypted_data_buf[1472] : encrypted_data_buf_next[1472];   // modexp_top.v(751)
    assign n8192 = rst ? encrypted_data_buf[1471] : encrypted_data_buf_next[1471];   // modexp_top.v(751)
    assign n8193 = rst ? encrypted_data_buf[1470] : encrypted_data_buf_next[1470];   // modexp_top.v(751)
    assign n8194 = rst ? encrypted_data_buf[1469] : encrypted_data_buf_next[1469];   // modexp_top.v(751)
    assign n8195 = rst ? encrypted_data_buf[1468] : encrypted_data_buf_next[1468];   // modexp_top.v(751)
    assign n8196 = rst ? encrypted_data_buf[1467] : encrypted_data_buf_next[1467];   // modexp_top.v(751)
    assign n8197 = rst ? encrypted_data_buf[1466] : encrypted_data_buf_next[1466];   // modexp_top.v(751)
    assign n8198 = rst ? encrypted_data_buf[1465] : encrypted_data_buf_next[1465];   // modexp_top.v(751)
    assign n8199 = rst ? encrypted_data_buf[1464] : encrypted_data_buf_next[1464];   // modexp_top.v(751)
    assign n8200 = rst ? encrypted_data_buf[1463] : encrypted_data_buf_next[1463];   // modexp_top.v(751)
    assign n8201 = rst ? encrypted_data_buf[1462] : encrypted_data_buf_next[1462];   // modexp_top.v(751)
    assign n8202 = rst ? encrypted_data_buf[1461] : encrypted_data_buf_next[1461];   // modexp_top.v(751)
    assign n8203 = rst ? encrypted_data_buf[1460] : encrypted_data_buf_next[1460];   // modexp_top.v(751)
    assign n8204 = rst ? encrypted_data_buf[1459] : encrypted_data_buf_next[1459];   // modexp_top.v(751)
    assign n8205 = rst ? encrypted_data_buf[1458] : encrypted_data_buf_next[1458];   // modexp_top.v(751)
    assign n8206 = rst ? encrypted_data_buf[1457] : encrypted_data_buf_next[1457];   // modexp_top.v(751)
    assign n8207 = rst ? encrypted_data_buf[1456] : encrypted_data_buf_next[1456];   // modexp_top.v(751)
    assign n8208 = rst ? encrypted_data_buf[1455] : encrypted_data_buf_next[1455];   // modexp_top.v(751)
    assign n8209 = rst ? encrypted_data_buf[1454] : encrypted_data_buf_next[1454];   // modexp_top.v(751)
    assign n8210 = rst ? encrypted_data_buf[1453] : encrypted_data_buf_next[1453];   // modexp_top.v(751)
    assign n8211 = rst ? encrypted_data_buf[1452] : encrypted_data_buf_next[1452];   // modexp_top.v(751)
    assign n8212 = rst ? encrypted_data_buf[1451] : encrypted_data_buf_next[1451];   // modexp_top.v(751)
    assign n8213 = rst ? encrypted_data_buf[1450] : encrypted_data_buf_next[1450];   // modexp_top.v(751)
    assign n8214 = rst ? encrypted_data_buf[1449] : encrypted_data_buf_next[1449];   // modexp_top.v(751)
    assign n8215 = rst ? encrypted_data_buf[1448] : encrypted_data_buf_next[1448];   // modexp_top.v(751)
    assign n8216 = rst ? encrypted_data_buf[1447] : encrypted_data_buf_next[1447];   // modexp_top.v(751)
    assign n8217 = rst ? encrypted_data_buf[1446] : encrypted_data_buf_next[1446];   // modexp_top.v(751)
    assign n8218 = rst ? encrypted_data_buf[1445] : encrypted_data_buf_next[1445];   // modexp_top.v(751)
    assign n8219 = rst ? encrypted_data_buf[1444] : encrypted_data_buf_next[1444];   // modexp_top.v(751)
    assign n8220 = rst ? encrypted_data_buf[1443] : encrypted_data_buf_next[1443];   // modexp_top.v(751)
    assign n8221 = rst ? encrypted_data_buf[1442] : encrypted_data_buf_next[1442];   // modexp_top.v(751)
    assign n8222 = rst ? encrypted_data_buf[1441] : encrypted_data_buf_next[1441];   // modexp_top.v(751)
    assign n8223 = rst ? encrypted_data_buf[1440] : encrypted_data_buf_next[1440];   // modexp_top.v(751)
    assign n8224 = rst ? encrypted_data_buf[1439] : encrypted_data_buf_next[1439];   // modexp_top.v(751)
    assign n8225 = rst ? encrypted_data_buf[1438] : encrypted_data_buf_next[1438];   // modexp_top.v(751)
    assign n8226 = rst ? encrypted_data_buf[1437] : encrypted_data_buf_next[1437];   // modexp_top.v(751)
    assign n8227 = rst ? encrypted_data_buf[1436] : encrypted_data_buf_next[1436];   // modexp_top.v(751)
    assign n8228 = rst ? encrypted_data_buf[1435] : encrypted_data_buf_next[1435];   // modexp_top.v(751)
    assign n8229 = rst ? encrypted_data_buf[1434] : encrypted_data_buf_next[1434];   // modexp_top.v(751)
    assign n8230 = rst ? encrypted_data_buf[1433] : encrypted_data_buf_next[1433];   // modexp_top.v(751)
    assign n8231 = rst ? encrypted_data_buf[1432] : encrypted_data_buf_next[1432];   // modexp_top.v(751)
    assign n8232 = rst ? encrypted_data_buf[1431] : encrypted_data_buf_next[1431];   // modexp_top.v(751)
    assign n8233 = rst ? encrypted_data_buf[1430] : encrypted_data_buf_next[1430];   // modexp_top.v(751)
    assign n8234 = rst ? encrypted_data_buf[1429] : encrypted_data_buf_next[1429];   // modexp_top.v(751)
    assign n8235 = rst ? encrypted_data_buf[1428] : encrypted_data_buf_next[1428];   // modexp_top.v(751)
    assign n8236 = rst ? encrypted_data_buf[1427] : encrypted_data_buf_next[1427];   // modexp_top.v(751)
    assign n8237 = rst ? encrypted_data_buf[1426] : encrypted_data_buf_next[1426];   // modexp_top.v(751)
    assign n8238 = rst ? encrypted_data_buf[1425] : encrypted_data_buf_next[1425];   // modexp_top.v(751)
    assign n8239 = rst ? encrypted_data_buf[1424] : encrypted_data_buf_next[1424];   // modexp_top.v(751)
    assign n8240 = rst ? encrypted_data_buf[1423] : encrypted_data_buf_next[1423];   // modexp_top.v(751)
    assign n8241 = rst ? encrypted_data_buf[1422] : encrypted_data_buf_next[1422];   // modexp_top.v(751)
    assign n8242 = rst ? encrypted_data_buf[1421] : encrypted_data_buf_next[1421];   // modexp_top.v(751)
    assign n8243 = rst ? encrypted_data_buf[1420] : encrypted_data_buf_next[1420];   // modexp_top.v(751)
    assign n8244 = rst ? encrypted_data_buf[1419] : encrypted_data_buf_next[1419];   // modexp_top.v(751)
    assign n8245 = rst ? encrypted_data_buf[1418] : encrypted_data_buf_next[1418];   // modexp_top.v(751)
    assign n8246 = rst ? encrypted_data_buf[1417] : encrypted_data_buf_next[1417];   // modexp_top.v(751)
    assign n8247 = rst ? encrypted_data_buf[1416] : encrypted_data_buf_next[1416];   // modexp_top.v(751)
    assign n8248 = rst ? encrypted_data_buf[1415] : encrypted_data_buf_next[1415];   // modexp_top.v(751)
    assign n8249 = rst ? encrypted_data_buf[1414] : encrypted_data_buf_next[1414];   // modexp_top.v(751)
    assign n8250 = rst ? encrypted_data_buf[1413] : encrypted_data_buf_next[1413];   // modexp_top.v(751)
    assign n8251 = rst ? encrypted_data_buf[1412] : encrypted_data_buf_next[1412];   // modexp_top.v(751)
    assign n8252 = rst ? encrypted_data_buf[1411] : encrypted_data_buf_next[1411];   // modexp_top.v(751)
    assign n8253 = rst ? encrypted_data_buf[1410] : encrypted_data_buf_next[1410];   // modexp_top.v(751)
    assign n8254 = rst ? encrypted_data_buf[1409] : encrypted_data_buf_next[1409];   // modexp_top.v(751)
    assign n8255 = rst ? encrypted_data_buf[1408] : encrypted_data_buf_next[1408];   // modexp_top.v(751)
    assign n8256 = rst ? encrypted_data_buf[1407] : encrypted_data_buf_next[1407];   // modexp_top.v(751)
    assign n8257 = rst ? encrypted_data_buf[1406] : encrypted_data_buf_next[1406];   // modexp_top.v(751)
    assign n8258 = rst ? encrypted_data_buf[1405] : encrypted_data_buf_next[1405];   // modexp_top.v(751)
    assign n8259 = rst ? encrypted_data_buf[1404] : encrypted_data_buf_next[1404];   // modexp_top.v(751)
    assign n8260 = rst ? encrypted_data_buf[1403] : encrypted_data_buf_next[1403];   // modexp_top.v(751)
    assign n8261 = rst ? encrypted_data_buf[1402] : encrypted_data_buf_next[1402];   // modexp_top.v(751)
    assign n8262 = rst ? encrypted_data_buf[1401] : encrypted_data_buf_next[1401];   // modexp_top.v(751)
    assign n8263 = rst ? encrypted_data_buf[1400] : encrypted_data_buf_next[1400];   // modexp_top.v(751)
    assign n8264 = rst ? encrypted_data_buf[1399] : encrypted_data_buf_next[1399];   // modexp_top.v(751)
    assign n8265 = rst ? encrypted_data_buf[1398] : encrypted_data_buf_next[1398];   // modexp_top.v(751)
    assign n8266 = rst ? encrypted_data_buf[1397] : encrypted_data_buf_next[1397];   // modexp_top.v(751)
    assign n8267 = rst ? encrypted_data_buf[1396] : encrypted_data_buf_next[1396];   // modexp_top.v(751)
    assign n8268 = rst ? encrypted_data_buf[1395] : encrypted_data_buf_next[1395];   // modexp_top.v(751)
    assign n8269 = rst ? encrypted_data_buf[1394] : encrypted_data_buf_next[1394];   // modexp_top.v(751)
    assign n8270 = rst ? encrypted_data_buf[1393] : encrypted_data_buf_next[1393];   // modexp_top.v(751)
    assign n8271 = rst ? encrypted_data_buf[1392] : encrypted_data_buf_next[1392];   // modexp_top.v(751)
    assign n8272 = rst ? encrypted_data_buf[1391] : encrypted_data_buf_next[1391];   // modexp_top.v(751)
    assign n8273 = rst ? encrypted_data_buf[1390] : encrypted_data_buf_next[1390];   // modexp_top.v(751)
    assign n8274 = rst ? encrypted_data_buf[1389] : encrypted_data_buf_next[1389];   // modexp_top.v(751)
    assign n8275 = rst ? encrypted_data_buf[1388] : encrypted_data_buf_next[1388];   // modexp_top.v(751)
    assign n8276 = rst ? encrypted_data_buf[1387] : encrypted_data_buf_next[1387];   // modexp_top.v(751)
    assign n8277 = rst ? encrypted_data_buf[1386] : encrypted_data_buf_next[1386];   // modexp_top.v(751)
    assign n8278 = rst ? encrypted_data_buf[1385] : encrypted_data_buf_next[1385];   // modexp_top.v(751)
    assign n8279 = rst ? encrypted_data_buf[1384] : encrypted_data_buf_next[1384];   // modexp_top.v(751)
    assign n8280 = rst ? encrypted_data_buf[1383] : encrypted_data_buf_next[1383];   // modexp_top.v(751)
    assign n8281 = rst ? encrypted_data_buf[1382] : encrypted_data_buf_next[1382];   // modexp_top.v(751)
    assign n8282 = rst ? encrypted_data_buf[1381] : encrypted_data_buf_next[1381];   // modexp_top.v(751)
    assign n8283 = rst ? encrypted_data_buf[1380] : encrypted_data_buf_next[1380];   // modexp_top.v(751)
    assign n8284 = rst ? encrypted_data_buf[1379] : encrypted_data_buf_next[1379];   // modexp_top.v(751)
    assign n8285 = rst ? encrypted_data_buf[1378] : encrypted_data_buf_next[1378];   // modexp_top.v(751)
    assign n8286 = rst ? encrypted_data_buf[1377] : encrypted_data_buf_next[1377];   // modexp_top.v(751)
    assign n8287 = rst ? encrypted_data_buf[1376] : encrypted_data_buf_next[1376];   // modexp_top.v(751)
    assign n8288 = rst ? encrypted_data_buf[1375] : encrypted_data_buf_next[1375];   // modexp_top.v(751)
    assign n8289 = rst ? encrypted_data_buf[1374] : encrypted_data_buf_next[1374];   // modexp_top.v(751)
    assign n8290 = rst ? encrypted_data_buf[1373] : encrypted_data_buf_next[1373];   // modexp_top.v(751)
    assign n8291 = rst ? encrypted_data_buf[1372] : encrypted_data_buf_next[1372];   // modexp_top.v(751)
    assign n8292 = rst ? encrypted_data_buf[1371] : encrypted_data_buf_next[1371];   // modexp_top.v(751)
    assign n8293 = rst ? encrypted_data_buf[1370] : encrypted_data_buf_next[1370];   // modexp_top.v(751)
    assign n8294 = rst ? encrypted_data_buf[1369] : encrypted_data_buf_next[1369];   // modexp_top.v(751)
    assign n8295 = rst ? encrypted_data_buf[1368] : encrypted_data_buf_next[1368];   // modexp_top.v(751)
    assign n8296 = rst ? encrypted_data_buf[1367] : encrypted_data_buf_next[1367];   // modexp_top.v(751)
    assign n8297 = rst ? encrypted_data_buf[1366] : encrypted_data_buf_next[1366];   // modexp_top.v(751)
    assign n8298 = rst ? encrypted_data_buf[1365] : encrypted_data_buf_next[1365];   // modexp_top.v(751)
    assign n8299 = rst ? encrypted_data_buf[1364] : encrypted_data_buf_next[1364];   // modexp_top.v(751)
    assign n8300 = rst ? encrypted_data_buf[1363] : encrypted_data_buf_next[1363];   // modexp_top.v(751)
    assign n8301 = rst ? encrypted_data_buf[1362] : encrypted_data_buf_next[1362];   // modexp_top.v(751)
    assign n8302 = rst ? encrypted_data_buf[1361] : encrypted_data_buf_next[1361];   // modexp_top.v(751)
    assign n8303 = rst ? encrypted_data_buf[1360] : encrypted_data_buf_next[1360];   // modexp_top.v(751)
    assign n8304 = rst ? encrypted_data_buf[1359] : encrypted_data_buf_next[1359];   // modexp_top.v(751)
    assign n8305 = rst ? encrypted_data_buf[1358] : encrypted_data_buf_next[1358];   // modexp_top.v(751)
    assign n8306 = rst ? encrypted_data_buf[1357] : encrypted_data_buf_next[1357];   // modexp_top.v(751)
    assign n8307 = rst ? encrypted_data_buf[1356] : encrypted_data_buf_next[1356];   // modexp_top.v(751)
    assign n8308 = rst ? encrypted_data_buf[1355] : encrypted_data_buf_next[1355];   // modexp_top.v(751)
    assign n8309 = rst ? encrypted_data_buf[1354] : encrypted_data_buf_next[1354];   // modexp_top.v(751)
    assign n8310 = rst ? encrypted_data_buf[1353] : encrypted_data_buf_next[1353];   // modexp_top.v(751)
    assign n8311 = rst ? encrypted_data_buf[1352] : encrypted_data_buf_next[1352];   // modexp_top.v(751)
    assign n8312 = rst ? encrypted_data_buf[1351] : encrypted_data_buf_next[1351];   // modexp_top.v(751)
    assign n8313 = rst ? encrypted_data_buf[1350] : encrypted_data_buf_next[1350];   // modexp_top.v(751)
    assign n8314 = rst ? encrypted_data_buf[1349] : encrypted_data_buf_next[1349];   // modexp_top.v(751)
    assign n8315 = rst ? encrypted_data_buf[1348] : encrypted_data_buf_next[1348];   // modexp_top.v(751)
    assign n8316 = rst ? encrypted_data_buf[1347] : encrypted_data_buf_next[1347];   // modexp_top.v(751)
    assign n8317 = rst ? encrypted_data_buf[1346] : encrypted_data_buf_next[1346];   // modexp_top.v(751)
    assign n8318 = rst ? encrypted_data_buf[1345] : encrypted_data_buf_next[1345];   // modexp_top.v(751)
    assign n8319 = rst ? encrypted_data_buf[1344] : encrypted_data_buf_next[1344];   // modexp_top.v(751)
    assign n8320 = rst ? encrypted_data_buf[1343] : encrypted_data_buf_next[1343];   // modexp_top.v(751)
    assign n8321 = rst ? encrypted_data_buf[1342] : encrypted_data_buf_next[1342];   // modexp_top.v(751)
    assign n8322 = rst ? encrypted_data_buf[1341] : encrypted_data_buf_next[1341];   // modexp_top.v(751)
    assign n8323 = rst ? encrypted_data_buf[1340] : encrypted_data_buf_next[1340];   // modexp_top.v(751)
    assign n8324 = rst ? encrypted_data_buf[1339] : encrypted_data_buf_next[1339];   // modexp_top.v(751)
    assign n8325 = rst ? encrypted_data_buf[1338] : encrypted_data_buf_next[1338];   // modexp_top.v(751)
    assign n8326 = rst ? encrypted_data_buf[1337] : encrypted_data_buf_next[1337];   // modexp_top.v(751)
    assign n8327 = rst ? encrypted_data_buf[1336] : encrypted_data_buf_next[1336];   // modexp_top.v(751)
    assign n8328 = rst ? encrypted_data_buf[1335] : encrypted_data_buf_next[1335];   // modexp_top.v(751)
    assign n8329 = rst ? encrypted_data_buf[1334] : encrypted_data_buf_next[1334];   // modexp_top.v(751)
    assign n8330 = rst ? encrypted_data_buf[1333] : encrypted_data_buf_next[1333];   // modexp_top.v(751)
    assign n8331 = rst ? encrypted_data_buf[1332] : encrypted_data_buf_next[1332];   // modexp_top.v(751)
    assign n8332 = rst ? encrypted_data_buf[1331] : encrypted_data_buf_next[1331];   // modexp_top.v(751)
    assign n8333 = rst ? encrypted_data_buf[1330] : encrypted_data_buf_next[1330];   // modexp_top.v(751)
    assign n8334 = rst ? encrypted_data_buf[1329] : encrypted_data_buf_next[1329];   // modexp_top.v(751)
    assign n8335 = rst ? encrypted_data_buf[1328] : encrypted_data_buf_next[1328];   // modexp_top.v(751)
    assign n8336 = rst ? encrypted_data_buf[1327] : encrypted_data_buf_next[1327];   // modexp_top.v(751)
    assign n8337 = rst ? encrypted_data_buf[1326] : encrypted_data_buf_next[1326];   // modexp_top.v(751)
    assign n8338 = rst ? encrypted_data_buf[1325] : encrypted_data_buf_next[1325];   // modexp_top.v(751)
    assign n8339 = rst ? encrypted_data_buf[1324] : encrypted_data_buf_next[1324];   // modexp_top.v(751)
    assign n8340 = rst ? encrypted_data_buf[1323] : encrypted_data_buf_next[1323];   // modexp_top.v(751)
    assign n8341 = rst ? encrypted_data_buf[1322] : encrypted_data_buf_next[1322];   // modexp_top.v(751)
    assign n8342 = rst ? encrypted_data_buf[1321] : encrypted_data_buf_next[1321];   // modexp_top.v(751)
    assign n8343 = rst ? encrypted_data_buf[1320] : encrypted_data_buf_next[1320];   // modexp_top.v(751)
    assign n8344 = rst ? encrypted_data_buf[1319] : encrypted_data_buf_next[1319];   // modexp_top.v(751)
    assign n8345 = rst ? encrypted_data_buf[1318] : encrypted_data_buf_next[1318];   // modexp_top.v(751)
    assign n8346 = rst ? encrypted_data_buf[1317] : encrypted_data_buf_next[1317];   // modexp_top.v(751)
    assign n8347 = rst ? encrypted_data_buf[1316] : encrypted_data_buf_next[1316];   // modexp_top.v(751)
    assign n8348 = rst ? encrypted_data_buf[1315] : encrypted_data_buf_next[1315];   // modexp_top.v(751)
    assign n8349 = rst ? encrypted_data_buf[1314] : encrypted_data_buf_next[1314];   // modexp_top.v(751)
    assign n8350 = rst ? encrypted_data_buf[1313] : encrypted_data_buf_next[1313];   // modexp_top.v(751)
    assign n8351 = rst ? encrypted_data_buf[1312] : encrypted_data_buf_next[1312];   // modexp_top.v(751)
    assign n8352 = rst ? encrypted_data_buf[1311] : encrypted_data_buf_next[1311];   // modexp_top.v(751)
    assign n8353 = rst ? encrypted_data_buf[1310] : encrypted_data_buf_next[1310];   // modexp_top.v(751)
    assign n8354 = rst ? encrypted_data_buf[1309] : encrypted_data_buf_next[1309];   // modexp_top.v(751)
    assign n8355 = rst ? encrypted_data_buf[1308] : encrypted_data_buf_next[1308];   // modexp_top.v(751)
    assign n8356 = rst ? encrypted_data_buf[1307] : encrypted_data_buf_next[1307];   // modexp_top.v(751)
    assign n8357 = rst ? encrypted_data_buf[1306] : encrypted_data_buf_next[1306];   // modexp_top.v(751)
    assign n8358 = rst ? encrypted_data_buf[1305] : encrypted_data_buf_next[1305];   // modexp_top.v(751)
    assign n8359 = rst ? encrypted_data_buf[1304] : encrypted_data_buf_next[1304];   // modexp_top.v(751)
    assign n8360 = rst ? encrypted_data_buf[1303] : encrypted_data_buf_next[1303];   // modexp_top.v(751)
    assign n8361 = rst ? encrypted_data_buf[1302] : encrypted_data_buf_next[1302];   // modexp_top.v(751)
    assign n8362 = rst ? encrypted_data_buf[1301] : encrypted_data_buf_next[1301];   // modexp_top.v(751)
    assign n8363 = rst ? encrypted_data_buf[1300] : encrypted_data_buf_next[1300];   // modexp_top.v(751)
    assign n8364 = rst ? encrypted_data_buf[1299] : encrypted_data_buf_next[1299];   // modexp_top.v(751)
    assign n8365 = rst ? encrypted_data_buf[1298] : encrypted_data_buf_next[1298];   // modexp_top.v(751)
    assign n8366 = rst ? encrypted_data_buf[1297] : encrypted_data_buf_next[1297];   // modexp_top.v(751)
    assign n8367 = rst ? encrypted_data_buf[1296] : encrypted_data_buf_next[1296];   // modexp_top.v(751)
    assign n8368 = rst ? encrypted_data_buf[1295] : encrypted_data_buf_next[1295];   // modexp_top.v(751)
    assign n8369 = rst ? encrypted_data_buf[1294] : encrypted_data_buf_next[1294];   // modexp_top.v(751)
    assign n8370 = rst ? encrypted_data_buf[1293] : encrypted_data_buf_next[1293];   // modexp_top.v(751)
    assign n8371 = rst ? encrypted_data_buf[1292] : encrypted_data_buf_next[1292];   // modexp_top.v(751)
    assign n8372 = rst ? encrypted_data_buf[1291] : encrypted_data_buf_next[1291];   // modexp_top.v(751)
    assign n8373 = rst ? encrypted_data_buf[1290] : encrypted_data_buf_next[1290];   // modexp_top.v(751)
    assign n8374 = rst ? encrypted_data_buf[1289] : encrypted_data_buf_next[1289];   // modexp_top.v(751)
    assign n8375 = rst ? encrypted_data_buf[1288] : encrypted_data_buf_next[1288];   // modexp_top.v(751)
    assign n8376 = rst ? encrypted_data_buf[1287] : encrypted_data_buf_next[1287];   // modexp_top.v(751)
    assign n8377 = rst ? encrypted_data_buf[1286] : encrypted_data_buf_next[1286];   // modexp_top.v(751)
    assign n8378 = rst ? encrypted_data_buf[1285] : encrypted_data_buf_next[1285];   // modexp_top.v(751)
    assign n8379 = rst ? encrypted_data_buf[1284] : encrypted_data_buf_next[1284];   // modexp_top.v(751)
    assign n8380 = rst ? encrypted_data_buf[1283] : encrypted_data_buf_next[1283];   // modexp_top.v(751)
    assign n8381 = rst ? encrypted_data_buf[1282] : encrypted_data_buf_next[1282];   // modexp_top.v(751)
    assign n8382 = rst ? encrypted_data_buf[1281] : encrypted_data_buf_next[1281];   // modexp_top.v(751)
    assign n8383 = rst ? encrypted_data_buf[1280] : encrypted_data_buf_next[1280];   // modexp_top.v(751)
    assign n8384 = rst ? encrypted_data_buf[1279] : encrypted_data_buf_next[1279];   // modexp_top.v(751)
    assign n8385 = rst ? encrypted_data_buf[1278] : encrypted_data_buf_next[1278];   // modexp_top.v(751)
    assign n8386 = rst ? encrypted_data_buf[1277] : encrypted_data_buf_next[1277];   // modexp_top.v(751)
    assign n8387 = rst ? encrypted_data_buf[1276] : encrypted_data_buf_next[1276];   // modexp_top.v(751)
    assign n8388 = rst ? encrypted_data_buf[1275] : encrypted_data_buf_next[1275];   // modexp_top.v(751)
    assign n8389 = rst ? encrypted_data_buf[1274] : encrypted_data_buf_next[1274];   // modexp_top.v(751)
    assign n8390 = rst ? encrypted_data_buf[1273] : encrypted_data_buf_next[1273];   // modexp_top.v(751)
    assign n8391 = rst ? encrypted_data_buf[1272] : encrypted_data_buf_next[1272];   // modexp_top.v(751)
    assign n8392 = rst ? encrypted_data_buf[1271] : encrypted_data_buf_next[1271];   // modexp_top.v(751)
    assign n8393 = rst ? encrypted_data_buf[1270] : encrypted_data_buf_next[1270];   // modexp_top.v(751)
    assign n8394 = rst ? encrypted_data_buf[1269] : encrypted_data_buf_next[1269];   // modexp_top.v(751)
    assign n8395 = rst ? encrypted_data_buf[1268] : encrypted_data_buf_next[1268];   // modexp_top.v(751)
    assign n8396 = rst ? encrypted_data_buf[1267] : encrypted_data_buf_next[1267];   // modexp_top.v(751)
    assign n8397 = rst ? encrypted_data_buf[1266] : encrypted_data_buf_next[1266];   // modexp_top.v(751)
    assign n8398 = rst ? encrypted_data_buf[1265] : encrypted_data_buf_next[1265];   // modexp_top.v(751)
    assign n8399 = rst ? encrypted_data_buf[1264] : encrypted_data_buf_next[1264];   // modexp_top.v(751)
    assign n8400 = rst ? encrypted_data_buf[1263] : encrypted_data_buf_next[1263];   // modexp_top.v(751)
    assign n8401 = rst ? encrypted_data_buf[1262] : encrypted_data_buf_next[1262];   // modexp_top.v(751)
    assign n8402 = rst ? encrypted_data_buf[1261] : encrypted_data_buf_next[1261];   // modexp_top.v(751)
    assign n8403 = rst ? encrypted_data_buf[1260] : encrypted_data_buf_next[1260];   // modexp_top.v(751)
    assign n8404 = rst ? encrypted_data_buf[1259] : encrypted_data_buf_next[1259];   // modexp_top.v(751)
    assign n8405 = rst ? encrypted_data_buf[1258] : encrypted_data_buf_next[1258];   // modexp_top.v(751)
    assign n8406 = rst ? encrypted_data_buf[1257] : encrypted_data_buf_next[1257];   // modexp_top.v(751)
    assign n8407 = rst ? encrypted_data_buf[1256] : encrypted_data_buf_next[1256];   // modexp_top.v(751)
    assign n8408 = rst ? encrypted_data_buf[1255] : encrypted_data_buf_next[1255];   // modexp_top.v(751)
    assign n8409 = rst ? encrypted_data_buf[1254] : encrypted_data_buf_next[1254];   // modexp_top.v(751)
    assign n8410 = rst ? encrypted_data_buf[1253] : encrypted_data_buf_next[1253];   // modexp_top.v(751)
    assign n8411 = rst ? encrypted_data_buf[1252] : encrypted_data_buf_next[1252];   // modexp_top.v(751)
    assign n8412 = rst ? encrypted_data_buf[1251] : encrypted_data_buf_next[1251];   // modexp_top.v(751)
    assign n8413 = rst ? encrypted_data_buf[1250] : encrypted_data_buf_next[1250];   // modexp_top.v(751)
    assign n8414 = rst ? encrypted_data_buf[1249] : encrypted_data_buf_next[1249];   // modexp_top.v(751)
    assign n8415 = rst ? encrypted_data_buf[1248] : encrypted_data_buf_next[1248];   // modexp_top.v(751)
    assign n8416 = rst ? encrypted_data_buf[1247] : encrypted_data_buf_next[1247];   // modexp_top.v(751)
    assign n8417 = rst ? encrypted_data_buf[1246] : encrypted_data_buf_next[1246];   // modexp_top.v(751)
    assign n8418 = rst ? encrypted_data_buf[1245] : encrypted_data_buf_next[1245];   // modexp_top.v(751)
    assign n8419 = rst ? encrypted_data_buf[1244] : encrypted_data_buf_next[1244];   // modexp_top.v(751)
    assign n8420 = rst ? encrypted_data_buf[1243] : encrypted_data_buf_next[1243];   // modexp_top.v(751)
    assign n8421 = rst ? encrypted_data_buf[1242] : encrypted_data_buf_next[1242];   // modexp_top.v(751)
    assign n8422 = rst ? encrypted_data_buf[1241] : encrypted_data_buf_next[1241];   // modexp_top.v(751)
    assign n8423 = rst ? encrypted_data_buf[1240] : encrypted_data_buf_next[1240];   // modexp_top.v(751)
    assign n8424 = rst ? encrypted_data_buf[1239] : encrypted_data_buf_next[1239];   // modexp_top.v(751)
    assign n8425 = rst ? encrypted_data_buf[1238] : encrypted_data_buf_next[1238];   // modexp_top.v(751)
    assign n8426 = rst ? encrypted_data_buf[1237] : encrypted_data_buf_next[1237];   // modexp_top.v(751)
    assign n8427 = rst ? encrypted_data_buf[1236] : encrypted_data_buf_next[1236];   // modexp_top.v(751)
    assign n8428 = rst ? encrypted_data_buf[1235] : encrypted_data_buf_next[1235];   // modexp_top.v(751)
    assign n8429 = rst ? encrypted_data_buf[1234] : encrypted_data_buf_next[1234];   // modexp_top.v(751)
    assign n8430 = rst ? encrypted_data_buf[1233] : encrypted_data_buf_next[1233];   // modexp_top.v(751)
    assign n8431 = rst ? encrypted_data_buf[1232] : encrypted_data_buf_next[1232];   // modexp_top.v(751)
    assign n8432 = rst ? encrypted_data_buf[1231] : encrypted_data_buf_next[1231];   // modexp_top.v(751)
    assign n8433 = rst ? encrypted_data_buf[1230] : encrypted_data_buf_next[1230];   // modexp_top.v(751)
    assign n8434 = rst ? encrypted_data_buf[1229] : encrypted_data_buf_next[1229];   // modexp_top.v(751)
    assign n8435 = rst ? encrypted_data_buf[1228] : encrypted_data_buf_next[1228];   // modexp_top.v(751)
    assign n8436 = rst ? encrypted_data_buf[1227] : encrypted_data_buf_next[1227];   // modexp_top.v(751)
    assign n8437 = rst ? encrypted_data_buf[1226] : encrypted_data_buf_next[1226];   // modexp_top.v(751)
    assign n8438 = rst ? encrypted_data_buf[1225] : encrypted_data_buf_next[1225];   // modexp_top.v(751)
    assign n8439 = rst ? encrypted_data_buf[1224] : encrypted_data_buf_next[1224];   // modexp_top.v(751)
    assign n8440 = rst ? encrypted_data_buf[1223] : encrypted_data_buf_next[1223];   // modexp_top.v(751)
    assign n8441 = rst ? encrypted_data_buf[1222] : encrypted_data_buf_next[1222];   // modexp_top.v(751)
    assign n8442 = rst ? encrypted_data_buf[1221] : encrypted_data_buf_next[1221];   // modexp_top.v(751)
    assign n8443 = rst ? encrypted_data_buf[1220] : encrypted_data_buf_next[1220];   // modexp_top.v(751)
    assign n8444 = rst ? encrypted_data_buf[1219] : encrypted_data_buf_next[1219];   // modexp_top.v(751)
    assign n8445 = rst ? encrypted_data_buf[1218] : encrypted_data_buf_next[1218];   // modexp_top.v(751)
    assign n8446 = rst ? encrypted_data_buf[1217] : encrypted_data_buf_next[1217];   // modexp_top.v(751)
    assign n8447 = rst ? encrypted_data_buf[1216] : encrypted_data_buf_next[1216];   // modexp_top.v(751)
    assign n8448 = rst ? encrypted_data_buf[1215] : encrypted_data_buf_next[1215];   // modexp_top.v(751)
    assign n8449 = rst ? encrypted_data_buf[1214] : encrypted_data_buf_next[1214];   // modexp_top.v(751)
    assign n8450 = rst ? encrypted_data_buf[1213] : encrypted_data_buf_next[1213];   // modexp_top.v(751)
    assign n8451 = rst ? encrypted_data_buf[1212] : encrypted_data_buf_next[1212];   // modexp_top.v(751)
    assign n8452 = rst ? encrypted_data_buf[1211] : encrypted_data_buf_next[1211];   // modexp_top.v(751)
    assign n8453 = rst ? encrypted_data_buf[1210] : encrypted_data_buf_next[1210];   // modexp_top.v(751)
    assign n8454 = rst ? encrypted_data_buf[1209] : encrypted_data_buf_next[1209];   // modexp_top.v(751)
    assign n8455 = rst ? encrypted_data_buf[1208] : encrypted_data_buf_next[1208];   // modexp_top.v(751)
    assign n8456 = rst ? encrypted_data_buf[1207] : encrypted_data_buf_next[1207];   // modexp_top.v(751)
    assign n8457 = rst ? encrypted_data_buf[1206] : encrypted_data_buf_next[1206];   // modexp_top.v(751)
    assign n8458 = rst ? encrypted_data_buf[1205] : encrypted_data_buf_next[1205];   // modexp_top.v(751)
    assign n8459 = rst ? encrypted_data_buf[1204] : encrypted_data_buf_next[1204];   // modexp_top.v(751)
    assign n8460 = rst ? encrypted_data_buf[1203] : encrypted_data_buf_next[1203];   // modexp_top.v(751)
    assign n8461 = rst ? encrypted_data_buf[1202] : encrypted_data_buf_next[1202];   // modexp_top.v(751)
    assign n8462 = rst ? encrypted_data_buf[1201] : encrypted_data_buf_next[1201];   // modexp_top.v(751)
    assign n8463 = rst ? encrypted_data_buf[1200] : encrypted_data_buf_next[1200];   // modexp_top.v(751)
    assign n8464 = rst ? encrypted_data_buf[1199] : encrypted_data_buf_next[1199];   // modexp_top.v(751)
    assign n8465 = rst ? encrypted_data_buf[1198] : encrypted_data_buf_next[1198];   // modexp_top.v(751)
    assign n8466 = rst ? encrypted_data_buf[1197] : encrypted_data_buf_next[1197];   // modexp_top.v(751)
    assign n8467 = rst ? encrypted_data_buf[1196] : encrypted_data_buf_next[1196];   // modexp_top.v(751)
    assign n8468 = rst ? encrypted_data_buf[1195] : encrypted_data_buf_next[1195];   // modexp_top.v(751)
    assign n8469 = rst ? encrypted_data_buf[1194] : encrypted_data_buf_next[1194];   // modexp_top.v(751)
    assign n8470 = rst ? encrypted_data_buf[1193] : encrypted_data_buf_next[1193];   // modexp_top.v(751)
    assign n8471 = rst ? encrypted_data_buf[1192] : encrypted_data_buf_next[1192];   // modexp_top.v(751)
    assign n8472 = rst ? encrypted_data_buf[1191] : encrypted_data_buf_next[1191];   // modexp_top.v(751)
    assign n8473 = rst ? encrypted_data_buf[1190] : encrypted_data_buf_next[1190];   // modexp_top.v(751)
    assign n8474 = rst ? encrypted_data_buf[1189] : encrypted_data_buf_next[1189];   // modexp_top.v(751)
    assign n8475 = rst ? encrypted_data_buf[1188] : encrypted_data_buf_next[1188];   // modexp_top.v(751)
    assign n8476 = rst ? encrypted_data_buf[1187] : encrypted_data_buf_next[1187];   // modexp_top.v(751)
    assign n8477 = rst ? encrypted_data_buf[1186] : encrypted_data_buf_next[1186];   // modexp_top.v(751)
    assign n8478 = rst ? encrypted_data_buf[1185] : encrypted_data_buf_next[1185];   // modexp_top.v(751)
    assign n8479 = rst ? encrypted_data_buf[1184] : encrypted_data_buf_next[1184];   // modexp_top.v(751)
    assign n8480 = rst ? encrypted_data_buf[1183] : encrypted_data_buf_next[1183];   // modexp_top.v(751)
    assign n8481 = rst ? encrypted_data_buf[1182] : encrypted_data_buf_next[1182];   // modexp_top.v(751)
    assign n8482 = rst ? encrypted_data_buf[1181] : encrypted_data_buf_next[1181];   // modexp_top.v(751)
    assign n8483 = rst ? encrypted_data_buf[1180] : encrypted_data_buf_next[1180];   // modexp_top.v(751)
    assign n8484 = rst ? encrypted_data_buf[1179] : encrypted_data_buf_next[1179];   // modexp_top.v(751)
    assign n8485 = rst ? encrypted_data_buf[1178] : encrypted_data_buf_next[1178];   // modexp_top.v(751)
    assign n8486 = rst ? encrypted_data_buf[1177] : encrypted_data_buf_next[1177];   // modexp_top.v(751)
    assign n8487 = rst ? encrypted_data_buf[1176] : encrypted_data_buf_next[1176];   // modexp_top.v(751)
    assign n8488 = rst ? encrypted_data_buf[1175] : encrypted_data_buf_next[1175];   // modexp_top.v(751)
    assign n8489 = rst ? encrypted_data_buf[1174] : encrypted_data_buf_next[1174];   // modexp_top.v(751)
    assign n8490 = rst ? encrypted_data_buf[1173] : encrypted_data_buf_next[1173];   // modexp_top.v(751)
    assign n8491 = rst ? encrypted_data_buf[1172] : encrypted_data_buf_next[1172];   // modexp_top.v(751)
    assign n8492 = rst ? encrypted_data_buf[1171] : encrypted_data_buf_next[1171];   // modexp_top.v(751)
    assign n8493 = rst ? encrypted_data_buf[1170] : encrypted_data_buf_next[1170];   // modexp_top.v(751)
    assign n8494 = rst ? encrypted_data_buf[1169] : encrypted_data_buf_next[1169];   // modexp_top.v(751)
    assign n8495 = rst ? encrypted_data_buf[1168] : encrypted_data_buf_next[1168];   // modexp_top.v(751)
    assign n8496 = rst ? encrypted_data_buf[1167] : encrypted_data_buf_next[1167];   // modexp_top.v(751)
    assign n8497 = rst ? encrypted_data_buf[1166] : encrypted_data_buf_next[1166];   // modexp_top.v(751)
    assign n8498 = rst ? encrypted_data_buf[1165] : encrypted_data_buf_next[1165];   // modexp_top.v(751)
    assign n8499 = rst ? encrypted_data_buf[1164] : encrypted_data_buf_next[1164];   // modexp_top.v(751)
    assign n8500 = rst ? encrypted_data_buf[1163] : encrypted_data_buf_next[1163];   // modexp_top.v(751)
    assign n8501 = rst ? encrypted_data_buf[1162] : encrypted_data_buf_next[1162];   // modexp_top.v(751)
    assign n8502 = rst ? encrypted_data_buf[1161] : encrypted_data_buf_next[1161];   // modexp_top.v(751)
    assign n8503 = rst ? encrypted_data_buf[1160] : encrypted_data_buf_next[1160];   // modexp_top.v(751)
    assign n8504 = rst ? encrypted_data_buf[1159] : encrypted_data_buf_next[1159];   // modexp_top.v(751)
    assign n8505 = rst ? encrypted_data_buf[1158] : encrypted_data_buf_next[1158];   // modexp_top.v(751)
    assign n8506 = rst ? encrypted_data_buf[1157] : encrypted_data_buf_next[1157];   // modexp_top.v(751)
    assign n8507 = rst ? encrypted_data_buf[1156] : encrypted_data_buf_next[1156];   // modexp_top.v(751)
    assign n8508 = rst ? encrypted_data_buf[1155] : encrypted_data_buf_next[1155];   // modexp_top.v(751)
    assign n8509 = rst ? encrypted_data_buf[1154] : encrypted_data_buf_next[1154];   // modexp_top.v(751)
    assign n8510 = rst ? encrypted_data_buf[1153] : encrypted_data_buf_next[1153];   // modexp_top.v(751)
    assign n8511 = rst ? encrypted_data_buf[1152] : encrypted_data_buf_next[1152];   // modexp_top.v(751)
    assign n8512 = rst ? encrypted_data_buf[1151] : encrypted_data_buf_next[1151];   // modexp_top.v(751)
    assign n8513 = rst ? encrypted_data_buf[1150] : encrypted_data_buf_next[1150];   // modexp_top.v(751)
    assign n8514 = rst ? encrypted_data_buf[1149] : encrypted_data_buf_next[1149];   // modexp_top.v(751)
    assign n8515 = rst ? encrypted_data_buf[1148] : encrypted_data_buf_next[1148];   // modexp_top.v(751)
    assign n8516 = rst ? encrypted_data_buf[1147] : encrypted_data_buf_next[1147];   // modexp_top.v(751)
    assign n8517 = rst ? encrypted_data_buf[1146] : encrypted_data_buf_next[1146];   // modexp_top.v(751)
    assign n8518 = rst ? encrypted_data_buf[1145] : encrypted_data_buf_next[1145];   // modexp_top.v(751)
    assign n8519 = rst ? encrypted_data_buf[1144] : encrypted_data_buf_next[1144];   // modexp_top.v(751)
    assign n8520 = rst ? encrypted_data_buf[1143] : encrypted_data_buf_next[1143];   // modexp_top.v(751)
    assign n8521 = rst ? encrypted_data_buf[1142] : encrypted_data_buf_next[1142];   // modexp_top.v(751)
    assign n8522 = rst ? encrypted_data_buf[1141] : encrypted_data_buf_next[1141];   // modexp_top.v(751)
    assign n8523 = rst ? encrypted_data_buf[1140] : encrypted_data_buf_next[1140];   // modexp_top.v(751)
    assign n8524 = rst ? encrypted_data_buf[1139] : encrypted_data_buf_next[1139];   // modexp_top.v(751)
    assign n8525 = rst ? encrypted_data_buf[1138] : encrypted_data_buf_next[1138];   // modexp_top.v(751)
    assign n8526 = rst ? encrypted_data_buf[1137] : encrypted_data_buf_next[1137];   // modexp_top.v(751)
    assign n8527 = rst ? encrypted_data_buf[1136] : encrypted_data_buf_next[1136];   // modexp_top.v(751)
    assign n8528 = rst ? encrypted_data_buf[1135] : encrypted_data_buf_next[1135];   // modexp_top.v(751)
    assign n8529 = rst ? encrypted_data_buf[1134] : encrypted_data_buf_next[1134];   // modexp_top.v(751)
    assign n8530 = rst ? encrypted_data_buf[1133] : encrypted_data_buf_next[1133];   // modexp_top.v(751)
    assign n8531 = rst ? encrypted_data_buf[1132] : encrypted_data_buf_next[1132];   // modexp_top.v(751)
    assign n8532 = rst ? encrypted_data_buf[1131] : encrypted_data_buf_next[1131];   // modexp_top.v(751)
    assign n8533 = rst ? encrypted_data_buf[1130] : encrypted_data_buf_next[1130];   // modexp_top.v(751)
    assign n8534 = rst ? encrypted_data_buf[1129] : encrypted_data_buf_next[1129];   // modexp_top.v(751)
    assign n8535 = rst ? encrypted_data_buf[1128] : encrypted_data_buf_next[1128];   // modexp_top.v(751)
    assign n8536 = rst ? encrypted_data_buf[1127] : encrypted_data_buf_next[1127];   // modexp_top.v(751)
    assign n8537 = rst ? encrypted_data_buf[1126] : encrypted_data_buf_next[1126];   // modexp_top.v(751)
    assign n8538 = rst ? encrypted_data_buf[1125] : encrypted_data_buf_next[1125];   // modexp_top.v(751)
    assign n8539 = rst ? encrypted_data_buf[1124] : encrypted_data_buf_next[1124];   // modexp_top.v(751)
    assign n8540 = rst ? encrypted_data_buf[1123] : encrypted_data_buf_next[1123];   // modexp_top.v(751)
    assign n8541 = rst ? encrypted_data_buf[1122] : encrypted_data_buf_next[1122];   // modexp_top.v(751)
    assign n8542 = rst ? encrypted_data_buf[1121] : encrypted_data_buf_next[1121];   // modexp_top.v(751)
    assign n8543 = rst ? encrypted_data_buf[1120] : encrypted_data_buf_next[1120];   // modexp_top.v(751)
    assign n8544 = rst ? encrypted_data_buf[1119] : encrypted_data_buf_next[1119];   // modexp_top.v(751)
    assign n8545 = rst ? encrypted_data_buf[1118] : encrypted_data_buf_next[1118];   // modexp_top.v(751)
    assign n8546 = rst ? encrypted_data_buf[1117] : encrypted_data_buf_next[1117];   // modexp_top.v(751)
    assign n8547 = rst ? encrypted_data_buf[1116] : encrypted_data_buf_next[1116];   // modexp_top.v(751)
    assign n8548 = rst ? encrypted_data_buf[1115] : encrypted_data_buf_next[1115];   // modexp_top.v(751)
    assign n8549 = rst ? encrypted_data_buf[1114] : encrypted_data_buf_next[1114];   // modexp_top.v(751)
    assign n8550 = rst ? encrypted_data_buf[1113] : encrypted_data_buf_next[1113];   // modexp_top.v(751)
    assign n8551 = rst ? encrypted_data_buf[1112] : encrypted_data_buf_next[1112];   // modexp_top.v(751)
    assign n8552 = rst ? encrypted_data_buf[1111] : encrypted_data_buf_next[1111];   // modexp_top.v(751)
    assign n8553 = rst ? encrypted_data_buf[1110] : encrypted_data_buf_next[1110];   // modexp_top.v(751)
    assign n8554 = rst ? encrypted_data_buf[1109] : encrypted_data_buf_next[1109];   // modexp_top.v(751)
    assign n8555 = rst ? encrypted_data_buf[1108] : encrypted_data_buf_next[1108];   // modexp_top.v(751)
    assign n8556 = rst ? encrypted_data_buf[1107] : encrypted_data_buf_next[1107];   // modexp_top.v(751)
    assign n8557 = rst ? encrypted_data_buf[1106] : encrypted_data_buf_next[1106];   // modexp_top.v(751)
    assign n8558 = rst ? encrypted_data_buf[1105] : encrypted_data_buf_next[1105];   // modexp_top.v(751)
    assign n8559 = rst ? encrypted_data_buf[1104] : encrypted_data_buf_next[1104];   // modexp_top.v(751)
    assign n8560 = rst ? encrypted_data_buf[1103] : encrypted_data_buf_next[1103];   // modexp_top.v(751)
    assign n8561 = rst ? encrypted_data_buf[1102] : encrypted_data_buf_next[1102];   // modexp_top.v(751)
    assign n8562 = rst ? encrypted_data_buf[1101] : encrypted_data_buf_next[1101];   // modexp_top.v(751)
    assign n8563 = rst ? encrypted_data_buf[1100] : encrypted_data_buf_next[1100];   // modexp_top.v(751)
    assign n8564 = rst ? encrypted_data_buf[1099] : encrypted_data_buf_next[1099];   // modexp_top.v(751)
    assign n8565 = rst ? encrypted_data_buf[1098] : encrypted_data_buf_next[1098];   // modexp_top.v(751)
    assign n8566 = rst ? encrypted_data_buf[1097] : encrypted_data_buf_next[1097];   // modexp_top.v(751)
    assign n8567 = rst ? encrypted_data_buf[1096] : encrypted_data_buf_next[1096];   // modexp_top.v(751)
    assign n8568 = rst ? encrypted_data_buf[1095] : encrypted_data_buf_next[1095];   // modexp_top.v(751)
    assign n8569 = rst ? encrypted_data_buf[1094] : encrypted_data_buf_next[1094];   // modexp_top.v(751)
    assign n8570 = rst ? encrypted_data_buf[1093] : encrypted_data_buf_next[1093];   // modexp_top.v(751)
    assign n8571 = rst ? encrypted_data_buf[1092] : encrypted_data_buf_next[1092];   // modexp_top.v(751)
    assign n8572 = rst ? encrypted_data_buf[1091] : encrypted_data_buf_next[1091];   // modexp_top.v(751)
    assign n8573 = rst ? encrypted_data_buf[1090] : encrypted_data_buf_next[1090];   // modexp_top.v(751)
    assign n8574 = rst ? encrypted_data_buf[1089] : encrypted_data_buf_next[1089];   // modexp_top.v(751)
    assign n8575 = rst ? encrypted_data_buf[1088] : encrypted_data_buf_next[1088];   // modexp_top.v(751)
    assign n8576 = rst ? encrypted_data_buf[1087] : encrypted_data_buf_next[1087];   // modexp_top.v(751)
    assign n8577 = rst ? encrypted_data_buf[1086] : encrypted_data_buf_next[1086];   // modexp_top.v(751)
    assign n8578 = rst ? encrypted_data_buf[1085] : encrypted_data_buf_next[1085];   // modexp_top.v(751)
    assign n8579 = rst ? encrypted_data_buf[1084] : encrypted_data_buf_next[1084];   // modexp_top.v(751)
    assign n8580 = rst ? encrypted_data_buf[1083] : encrypted_data_buf_next[1083];   // modexp_top.v(751)
    assign n8581 = rst ? encrypted_data_buf[1082] : encrypted_data_buf_next[1082];   // modexp_top.v(751)
    assign n8582 = rst ? encrypted_data_buf[1081] : encrypted_data_buf_next[1081];   // modexp_top.v(751)
    assign n8583 = rst ? encrypted_data_buf[1080] : encrypted_data_buf_next[1080];   // modexp_top.v(751)
    assign n8584 = rst ? encrypted_data_buf[1079] : encrypted_data_buf_next[1079];   // modexp_top.v(751)
    assign n8585 = rst ? encrypted_data_buf[1078] : encrypted_data_buf_next[1078];   // modexp_top.v(751)
    assign n8586 = rst ? encrypted_data_buf[1077] : encrypted_data_buf_next[1077];   // modexp_top.v(751)
    assign n8587 = rst ? encrypted_data_buf[1076] : encrypted_data_buf_next[1076];   // modexp_top.v(751)
    assign n8588 = rst ? encrypted_data_buf[1075] : encrypted_data_buf_next[1075];   // modexp_top.v(751)
    assign n8589 = rst ? encrypted_data_buf[1074] : encrypted_data_buf_next[1074];   // modexp_top.v(751)
    assign n8590 = rst ? encrypted_data_buf[1073] : encrypted_data_buf_next[1073];   // modexp_top.v(751)
    assign n8591 = rst ? encrypted_data_buf[1072] : encrypted_data_buf_next[1072];   // modexp_top.v(751)
    assign n8592 = rst ? encrypted_data_buf[1071] : encrypted_data_buf_next[1071];   // modexp_top.v(751)
    assign n8593 = rst ? encrypted_data_buf[1070] : encrypted_data_buf_next[1070];   // modexp_top.v(751)
    assign n8594 = rst ? encrypted_data_buf[1069] : encrypted_data_buf_next[1069];   // modexp_top.v(751)
    assign n8595 = rst ? encrypted_data_buf[1068] : encrypted_data_buf_next[1068];   // modexp_top.v(751)
    assign n8596 = rst ? encrypted_data_buf[1067] : encrypted_data_buf_next[1067];   // modexp_top.v(751)
    assign n8597 = rst ? encrypted_data_buf[1066] : encrypted_data_buf_next[1066];   // modexp_top.v(751)
    assign n8598 = rst ? encrypted_data_buf[1065] : encrypted_data_buf_next[1065];   // modexp_top.v(751)
    assign n8599 = rst ? encrypted_data_buf[1064] : encrypted_data_buf_next[1064];   // modexp_top.v(751)
    assign n8600 = rst ? encrypted_data_buf[1063] : encrypted_data_buf_next[1063];   // modexp_top.v(751)
    assign n8601 = rst ? encrypted_data_buf[1062] : encrypted_data_buf_next[1062];   // modexp_top.v(751)
    assign n8602 = rst ? encrypted_data_buf[1061] : encrypted_data_buf_next[1061];   // modexp_top.v(751)
    assign n8603 = rst ? encrypted_data_buf[1060] : encrypted_data_buf_next[1060];   // modexp_top.v(751)
    assign n8604 = rst ? encrypted_data_buf[1059] : encrypted_data_buf_next[1059];   // modexp_top.v(751)
    assign n8605 = rst ? encrypted_data_buf[1058] : encrypted_data_buf_next[1058];   // modexp_top.v(751)
    assign n8606 = rst ? encrypted_data_buf[1057] : encrypted_data_buf_next[1057];   // modexp_top.v(751)
    assign n8607 = rst ? encrypted_data_buf[1056] : encrypted_data_buf_next[1056];   // modexp_top.v(751)
    assign n8608 = rst ? encrypted_data_buf[1055] : encrypted_data_buf_next[1055];   // modexp_top.v(751)
    assign n8609 = rst ? encrypted_data_buf[1054] : encrypted_data_buf_next[1054];   // modexp_top.v(751)
    assign n8610 = rst ? encrypted_data_buf[1053] : encrypted_data_buf_next[1053];   // modexp_top.v(751)
    assign n8611 = rst ? encrypted_data_buf[1052] : encrypted_data_buf_next[1052];   // modexp_top.v(751)
    assign n8612 = rst ? encrypted_data_buf[1051] : encrypted_data_buf_next[1051];   // modexp_top.v(751)
    assign n8613 = rst ? encrypted_data_buf[1050] : encrypted_data_buf_next[1050];   // modexp_top.v(751)
    assign n8614 = rst ? encrypted_data_buf[1049] : encrypted_data_buf_next[1049];   // modexp_top.v(751)
    assign n8615 = rst ? encrypted_data_buf[1048] : encrypted_data_buf_next[1048];   // modexp_top.v(751)
    assign n8616 = rst ? encrypted_data_buf[1047] : encrypted_data_buf_next[1047];   // modexp_top.v(751)
    assign n8617 = rst ? encrypted_data_buf[1046] : encrypted_data_buf_next[1046];   // modexp_top.v(751)
    assign n8618 = rst ? encrypted_data_buf[1045] : encrypted_data_buf_next[1045];   // modexp_top.v(751)
    assign n8619 = rst ? encrypted_data_buf[1044] : encrypted_data_buf_next[1044];   // modexp_top.v(751)
    assign n8620 = rst ? encrypted_data_buf[1043] : encrypted_data_buf_next[1043];   // modexp_top.v(751)
    assign n8621 = rst ? encrypted_data_buf[1042] : encrypted_data_buf_next[1042];   // modexp_top.v(751)
    assign n8622 = rst ? encrypted_data_buf[1041] : encrypted_data_buf_next[1041];   // modexp_top.v(751)
    assign n8623 = rst ? encrypted_data_buf[1040] : encrypted_data_buf_next[1040];   // modexp_top.v(751)
    assign n8624 = rst ? encrypted_data_buf[1039] : encrypted_data_buf_next[1039];   // modexp_top.v(751)
    assign n8625 = rst ? encrypted_data_buf[1038] : encrypted_data_buf_next[1038];   // modexp_top.v(751)
    assign n8626 = rst ? encrypted_data_buf[1037] : encrypted_data_buf_next[1037];   // modexp_top.v(751)
    assign n8627 = rst ? encrypted_data_buf[1036] : encrypted_data_buf_next[1036];   // modexp_top.v(751)
    assign n8628 = rst ? encrypted_data_buf[1035] : encrypted_data_buf_next[1035];   // modexp_top.v(751)
    assign n8629 = rst ? encrypted_data_buf[1034] : encrypted_data_buf_next[1034];   // modexp_top.v(751)
    assign n8630 = rst ? encrypted_data_buf[1033] : encrypted_data_buf_next[1033];   // modexp_top.v(751)
    assign n8631 = rst ? encrypted_data_buf[1032] : encrypted_data_buf_next[1032];   // modexp_top.v(751)
    assign n8632 = rst ? encrypted_data_buf[1031] : encrypted_data_buf_next[1031];   // modexp_top.v(751)
    assign n8633 = rst ? encrypted_data_buf[1030] : encrypted_data_buf_next[1030];   // modexp_top.v(751)
    assign n8634 = rst ? encrypted_data_buf[1029] : encrypted_data_buf_next[1029];   // modexp_top.v(751)
    assign n8635 = rst ? encrypted_data_buf[1028] : encrypted_data_buf_next[1028];   // modexp_top.v(751)
    assign n8636 = rst ? encrypted_data_buf[1027] : encrypted_data_buf_next[1027];   // modexp_top.v(751)
    assign n8637 = rst ? encrypted_data_buf[1026] : encrypted_data_buf_next[1026];   // modexp_top.v(751)
    assign n8638 = rst ? encrypted_data_buf[1025] : encrypted_data_buf_next[1025];   // modexp_top.v(751)
    assign n8639 = rst ? encrypted_data_buf[1024] : encrypted_data_buf_next[1024];   // modexp_top.v(751)
    assign n8640 = rst ? encrypted_data_buf[1023] : encrypted_data_buf_next[1023];   // modexp_top.v(751)
    assign n8641 = rst ? encrypted_data_buf[1022] : encrypted_data_buf_next[1022];   // modexp_top.v(751)
    assign n8642 = rst ? encrypted_data_buf[1021] : encrypted_data_buf_next[1021];   // modexp_top.v(751)
    assign n8643 = rst ? encrypted_data_buf[1020] : encrypted_data_buf_next[1020];   // modexp_top.v(751)
    assign n8644 = rst ? encrypted_data_buf[1019] : encrypted_data_buf_next[1019];   // modexp_top.v(751)
    assign n8645 = rst ? encrypted_data_buf[1018] : encrypted_data_buf_next[1018];   // modexp_top.v(751)
    assign n8646 = rst ? encrypted_data_buf[1017] : encrypted_data_buf_next[1017];   // modexp_top.v(751)
    assign n8647 = rst ? encrypted_data_buf[1016] : encrypted_data_buf_next[1016];   // modexp_top.v(751)
    assign n8648 = rst ? encrypted_data_buf[1015] : encrypted_data_buf_next[1015];   // modexp_top.v(751)
    assign n8649 = rst ? encrypted_data_buf[1014] : encrypted_data_buf_next[1014];   // modexp_top.v(751)
    assign n8650 = rst ? encrypted_data_buf[1013] : encrypted_data_buf_next[1013];   // modexp_top.v(751)
    assign n8651 = rst ? encrypted_data_buf[1012] : encrypted_data_buf_next[1012];   // modexp_top.v(751)
    assign n8652 = rst ? encrypted_data_buf[1011] : encrypted_data_buf_next[1011];   // modexp_top.v(751)
    assign n8653 = rst ? encrypted_data_buf[1010] : encrypted_data_buf_next[1010];   // modexp_top.v(751)
    assign n8654 = rst ? encrypted_data_buf[1009] : encrypted_data_buf_next[1009];   // modexp_top.v(751)
    assign n8655 = rst ? encrypted_data_buf[1008] : encrypted_data_buf_next[1008];   // modexp_top.v(751)
    assign n8656 = rst ? encrypted_data_buf[1007] : encrypted_data_buf_next[1007];   // modexp_top.v(751)
    assign n8657 = rst ? encrypted_data_buf[1006] : encrypted_data_buf_next[1006];   // modexp_top.v(751)
    assign n8658 = rst ? encrypted_data_buf[1005] : encrypted_data_buf_next[1005];   // modexp_top.v(751)
    assign n8659 = rst ? encrypted_data_buf[1004] : encrypted_data_buf_next[1004];   // modexp_top.v(751)
    assign n8660 = rst ? encrypted_data_buf[1003] : encrypted_data_buf_next[1003];   // modexp_top.v(751)
    assign n8661 = rst ? encrypted_data_buf[1002] : encrypted_data_buf_next[1002];   // modexp_top.v(751)
    assign n8662 = rst ? encrypted_data_buf[1001] : encrypted_data_buf_next[1001];   // modexp_top.v(751)
    assign n8663 = rst ? encrypted_data_buf[1000] : encrypted_data_buf_next[1000];   // modexp_top.v(751)
    assign n8664 = rst ? encrypted_data_buf[999] : encrypted_data_buf_next[999];   // modexp_top.v(751)
    assign n8665 = rst ? encrypted_data_buf[998] : encrypted_data_buf_next[998];   // modexp_top.v(751)
    assign n8666 = rst ? encrypted_data_buf[997] : encrypted_data_buf_next[997];   // modexp_top.v(751)
    assign n8667 = rst ? encrypted_data_buf[996] : encrypted_data_buf_next[996];   // modexp_top.v(751)
    assign n8668 = rst ? encrypted_data_buf[995] : encrypted_data_buf_next[995];   // modexp_top.v(751)
    assign n8669 = rst ? encrypted_data_buf[994] : encrypted_data_buf_next[994];   // modexp_top.v(751)
    assign n8670 = rst ? encrypted_data_buf[993] : encrypted_data_buf_next[993];   // modexp_top.v(751)
    assign n8671 = rst ? encrypted_data_buf[992] : encrypted_data_buf_next[992];   // modexp_top.v(751)
    assign n8672 = rst ? encrypted_data_buf[991] : encrypted_data_buf_next[991];   // modexp_top.v(751)
    assign n8673 = rst ? encrypted_data_buf[990] : encrypted_data_buf_next[990];   // modexp_top.v(751)
    assign n8674 = rst ? encrypted_data_buf[989] : encrypted_data_buf_next[989];   // modexp_top.v(751)
    assign n8675 = rst ? encrypted_data_buf[988] : encrypted_data_buf_next[988];   // modexp_top.v(751)
    assign n8676 = rst ? encrypted_data_buf[987] : encrypted_data_buf_next[987];   // modexp_top.v(751)
    assign n8677 = rst ? encrypted_data_buf[986] : encrypted_data_buf_next[986];   // modexp_top.v(751)
    assign n8678 = rst ? encrypted_data_buf[985] : encrypted_data_buf_next[985];   // modexp_top.v(751)
    assign n8679 = rst ? encrypted_data_buf[984] : encrypted_data_buf_next[984];   // modexp_top.v(751)
    assign n8680 = rst ? encrypted_data_buf[983] : encrypted_data_buf_next[983];   // modexp_top.v(751)
    assign n8681 = rst ? encrypted_data_buf[982] : encrypted_data_buf_next[982];   // modexp_top.v(751)
    assign n8682 = rst ? encrypted_data_buf[981] : encrypted_data_buf_next[981];   // modexp_top.v(751)
    assign n8683 = rst ? encrypted_data_buf[980] : encrypted_data_buf_next[980];   // modexp_top.v(751)
    assign n8684 = rst ? encrypted_data_buf[979] : encrypted_data_buf_next[979];   // modexp_top.v(751)
    assign n8685 = rst ? encrypted_data_buf[978] : encrypted_data_buf_next[978];   // modexp_top.v(751)
    assign n8686 = rst ? encrypted_data_buf[977] : encrypted_data_buf_next[977];   // modexp_top.v(751)
    assign n8687 = rst ? encrypted_data_buf[976] : encrypted_data_buf_next[976];   // modexp_top.v(751)
    assign n8688 = rst ? encrypted_data_buf[975] : encrypted_data_buf_next[975];   // modexp_top.v(751)
    assign n8689 = rst ? encrypted_data_buf[974] : encrypted_data_buf_next[974];   // modexp_top.v(751)
    assign n8690 = rst ? encrypted_data_buf[973] : encrypted_data_buf_next[973];   // modexp_top.v(751)
    assign n8691 = rst ? encrypted_data_buf[972] : encrypted_data_buf_next[972];   // modexp_top.v(751)
    assign n8692 = rst ? encrypted_data_buf[971] : encrypted_data_buf_next[971];   // modexp_top.v(751)
    assign n8693 = rst ? encrypted_data_buf[970] : encrypted_data_buf_next[970];   // modexp_top.v(751)
    assign n8694 = rst ? encrypted_data_buf[969] : encrypted_data_buf_next[969];   // modexp_top.v(751)
    assign n8695 = rst ? encrypted_data_buf[968] : encrypted_data_buf_next[968];   // modexp_top.v(751)
    assign n8696 = rst ? encrypted_data_buf[967] : encrypted_data_buf_next[967];   // modexp_top.v(751)
    assign n8697 = rst ? encrypted_data_buf[966] : encrypted_data_buf_next[966];   // modexp_top.v(751)
    assign n8698 = rst ? encrypted_data_buf[965] : encrypted_data_buf_next[965];   // modexp_top.v(751)
    assign n8699 = rst ? encrypted_data_buf[964] : encrypted_data_buf_next[964];   // modexp_top.v(751)
    assign n8700 = rst ? encrypted_data_buf[963] : encrypted_data_buf_next[963];   // modexp_top.v(751)
    assign n8701 = rst ? encrypted_data_buf[962] : encrypted_data_buf_next[962];   // modexp_top.v(751)
    assign n8702 = rst ? encrypted_data_buf[961] : encrypted_data_buf_next[961];   // modexp_top.v(751)
    assign n8703 = rst ? encrypted_data_buf[960] : encrypted_data_buf_next[960];   // modexp_top.v(751)
    assign n8704 = rst ? encrypted_data_buf[959] : encrypted_data_buf_next[959];   // modexp_top.v(751)
    assign n8705 = rst ? encrypted_data_buf[958] : encrypted_data_buf_next[958];   // modexp_top.v(751)
    assign n8706 = rst ? encrypted_data_buf[957] : encrypted_data_buf_next[957];   // modexp_top.v(751)
    assign n8707 = rst ? encrypted_data_buf[956] : encrypted_data_buf_next[956];   // modexp_top.v(751)
    assign n8708 = rst ? encrypted_data_buf[955] : encrypted_data_buf_next[955];   // modexp_top.v(751)
    assign n8709 = rst ? encrypted_data_buf[954] : encrypted_data_buf_next[954];   // modexp_top.v(751)
    assign n8710 = rst ? encrypted_data_buf[953] : encrypted_data_buf_next[953];   // modexp_top.v(751)
    assign n8711 = rst ? encrypted_data_buf[952] : encrypted_data_buf_next[952];   // modexp_top.v(751)
    assign n8712 = rst ? encrypted_data_buf[951] : encrypted_data_buf_next[951];   // modexp_top.v(751)
    assign n8713 = rst ? encrypted_data_buf[950] : encrypted_data_buf_next[950];   // modexp_top.v(751)
    assign n8714 = rst ? encrypted_data_buf[949] : encrypted_data_buf_next[949];   // modexp_top.v(751)
    assign n8715 = rst ? encrypted_data_buf[948] : encrypted_data_buf_next[948];   // modexp_top.v(751)
    assign n8716 = rst ? encrypted_data_buf[947] : encrypted_data_buf_next[947];   // modexp_top.v(751)
    assign n8717 = rst ? encrypted_data_buf[946] : encrypted_data_buf_next[946];   // modexp_top.v(751)
    assign n8718 = rst ? encrypted_data_buf[945] : encrypted_data_buf_next[945];   // modexp_top.v(751)
    assign n8719 = rst ? encrypted_data_buf[944] : encrypted_data_buf_next[944];   // modexp_top.v(751)
    assign n8720 = rst ? encrypted_data_buf[943] : encrypted_data_buf_next[943];   // modexp_top.v(751)
    assign n8721 = rst ? encrypted_data_buf[942] : encrypted_data_buf_next[942];   // modexp_top.v(751)
    assign n8722 = rst ? encrypted_data_buf[941] : encrypted_data_buf_next[941];   // modexp_top.v(751)
    assign n8723 = rst ? encrypted_data_buf[940] : encrypted_data_buf_next[940];   // modexp_top.v(751)
    assign n8724 = rst ? encrypted_data_buf[939] : encrypted_data_buf_next[939];   // modexp_top.v(751)
    assign n8725 = rst ? encrypted_data_buf[938] : encrypted_data_buf_next[938];   // modexp_top.v(751)
    assign n8726 = rst ? encrypted_data_buf[937] : encrypted_data_buf_next[937];   // modexp_top.v(751)
    assign n8727 = rst ? encrypted_data_buf[936] : encrypted_data_buf_next[936];   // modexp_top.v(751)
    assign n8728 = rst ? encrypted_data_buf[935] : encrypted_data_buf_next[935];   // modexp_top.v(751)
    assign n8729 = rst ? encrypted_data_buf[934] : encrypted_data_buf_next[934];   // modexp_top.v(751)
    assign n8730 = rst ? encrypted_data_buf[933] : encrypted_data_buf_next[933];   // modexp_top.v(751)
    assign n8731 = rst ? encrypted_data_buf[932] : encrypted_data_buf_next[932];   // modexp_top.v(751)
    assign n8732 = rst ? encrypted_data_buf[931] : encrypted_data_buf_next[931];   // modexp_top.v(751)
    assign n8733 = rst ? encrypted_data_buf[930] : encrypted_data_buf_next[930];   // modexp_top.v(751)
    assign n8734 = rst ? encrypted_data_buf[929] : encrypted_data_buf_next[929];   // modexp_top.v(751)
    assign n8735 = rst ? encrypted_data_buf[928] : encrypted_data_buf_next[928];   // modexp_top.v(751)
    assign n8736 = rst ? encrypted_data_buf[927] : encrypted_data_buf_next[927];   // modexp_top.v(751)
    assign n8737 = rst ? encrypted_data_buf[926] : encrypted_data_buf_next[926];   // modexp_top.v(751)
    assign n8738 = rst ? encrypted_data_buf[925] : encrypted_data_buf_next[925];   // modexp_top.v(751)
    assign n8739 = rst ? encrypted_data_buf[924] : encrypted_data_buf_next[924];   // modexp_top.v(751)
    assign n8740 = rst ? encrypted_data_buf[923] : encrypted_data_buf_next[923];   // modexp_top.v(751)
    assign n8741 = rst ? encrypted_data_buf[922] : encrypted_data_buf_next[922];   // modexp_top.v(751)
    assign n8742 = rst ? encrypted_data_buf[921] : encrypted_data_buf_next[921];   // modexp_top.v(751)
    assign n8743 = rst ? encrypted_data_buf[920] : encrypted_data_buf_next[920];   // modexp_top.v(751)
    assign n8744 = rst ? encrypted_data_buf[919] : encrypted_data_buf_next[919];   // modexp_top.v(751)
    assign n8745 = rst ? encrypted_data_buf[918] : encrypted_data_buf_next[918];   // modexp_top.v(751)
    assign n8746 = rst ? encrypted_data_buf[917] : encrypted_data_buf_next[917];   // modexp_top.v(751)
    assign n8747 = rst ? encrypted_data_buf[916] : encrypted_data_buf_next[916];   // modexp_top.v(751)
    assign n8748 = rst ? encrypted_data_buf[915] : encrypted_data_buf_next[915];   // modexp_top.v(751)
    assign n8749 = rst ? encrypted_data_buf[914] : encrypted_data_buf_next[914];   // modexp_top.v(751)
    assign n8750 = rst ? encrypted_data_buf[913] : encrypted_data_buf_next[913];   // modexp_top.v(751)
    assign n8751 = rst ? encrypted_data_buf[912] : encrypted_data_buf_next[912];   // modexp_top.v(751)
    assign n8752 = rst ? encrypted_data_buf[911] : encrypted_data_buf_next[911];   // modexp_top.v(751)
    assign n8753 = rst ? encrypted_data_buf[910] : encrypted_data_buf_next[910];   // modexp_top.v(751)
    assign n8754 = rst ? encrypted_data_buf[909] : encrypted_data_buf_next[909];   // modexp_top.v(751)
    assign n8755 = rst ? encrypted_data_buf[908] : encrypted_data_buf_next[908];   // modexp_top.v(751)
    assign n8756 = rst ? encrypted_data_buf[907] : encrypted_data_buf_next[907];   // modexp_top.v(751)
    assign n8757 = rst ? encrypted_data_buf[906] : encrypted_data_buf_next[906];   // modexp_top.v(751)
    assign n8758 = rst ? encrypted_data_buf[905] : encrypted_data_buf_next[905];   // modexp_top.v(751)
    assign n8759 = rst ? encrypted_data_buf[904] : encrypted_data_buf_next[904];   // modexp_top.v(751)
    assign n8760 = rst ? encrypted_data_buf[903] : encrypted_data_buf_next[903];   // modexp_top.v(751)
    assign n8761 = rst ? encrypted_data_buf[902] : encrypted_data_buf_next[902];   // modexp_top.v(751)
    assign n8762 = rst ? encrypted_data_buf[901] : encrypted_data_buf_next[901];   // modexp_top.v(751)
    assign n8763 = rst ? encrypted_data_buf[900] : encrypted_data_buf_next[900];   // modexp_top.v(751)
    assign n8764 = rst ? encrypted_data_buf[899] : encrypted_data_buf_next[899];   // modexp_top.v(751)
    assign n8765 = rst ? encrypted_data_buf[898] : encrypted_data_buf_next[898];   // modexp_top.v(751)
    assign n8766 = rst ? encrypted_data_buf[897] : encrypted_data_buf_next[897];   // modexp_top.v(751)
    assign n8767 = rst ? encrypted_data_buf[896] : encrypted_data_buf_next[896];   // modexp_top.v(751)
    assign n8768 = rst ? encrypted_data_buf[895] : encrypted_data_buf_next[895];   // modexp_top.v(751)
    assign n8769 = rst ? encrypted_data_buf[894] : encrypted_data_buf_next[894];   // modexp_top.v(751)
    assign n8770 = rst ? encrypted_data_buf[893] : encrypted_data_buf_next[893];   // modexp_top.v(751)
    assign n8771 = rst ? encrypted_data_buf[892] : encrypted_data_buf_next[892];   // modexp_top.v(751)
    assign n8772 = rst ? encrypted_data_buf[891] : encrypted_data_buf_next[891];   // modexp_top.v(751)
    assign n8773 = rst ? encrypted_data_buf[890] : encrypted_data_buf_next[890];   // modexp_top.v(751)
    assign n8774 = rst ? encrypted_data_buf[889] : encrypted_data_buf_next[889];   // modexp_top.v(751)
    assign n8775 = rst ? encrypted_data_buf[888] : encrypted_data_buf_next[888];   // modexp_top.v(751)
    assign n8776 = rst ? encrypted_data_buf[887] : encrypted_data_buf_next[887];   // modexp_top.v(751)
    assign n8777 = rst ? encrypted_data_buf[886] : encrypted_data_buf_next[886];   // modexp_top.v(751)
    assign n8778 = rst ? encrypted_data_buf[885] : encrypted_data_buf_next[885];   // modexp_top.v(751)
    assign n8779 = rst ? encrypted_data_buf[884] : encrypted_data_buf_next[884];   // modexp_top.v(751)
    assign n8780 = rst ? encrypted_data_buf[883] : encrypted_data_buf_next[883];   // modexp_top.v(751)
    assign n8781 = rst ? encrypted_data_buf[882] : encrypted_data_buf_next[882];   // modexp_top.v(751)
    assign n8782 = rst ? encrypted_data_buf[881] : encrypted_data_buf_next[881];   // modexp_top.v(751)
    assign n8783 = rst ? encrypted_data_buf[880] : encrypted_data_buf_next[880];   // modexp_top.v(751)
    assign n8784 = rst ? encrypted_data_buf[879] : encrypted_data_buf_next[879];   // modexp_top.v(751)
    assign n8785 = rst ? encrypted_data_buf[878] : encrypted_data_buf_next[878];   // modexp_top.v(751)
    assign n8786 = rst ? encrypted_data_buf[877] : encrypted_data_buf_next[877];   // modexp_top.v(751)
    assign n8787 = rst ? encrypted_data_buf[876] : encrypted_data_buf_next[876];   // modexp_top.v(751)
    assign n8788 = rst ? encrypted_data_buf[875] : encrypted_data_buf_next[875];   // modexp_top.v(751)
    assign n8789 = rst ? encrypted_data_buf[874] : encrypted_data_buf_next[874];   // modexp_top.v(751)
    assign n8790 = rst ? encrypted_data_buf[873] : encrypted_data_buf_next[873];   // modexp_top.v(751)
    assign n8791 = rst ? encrypted_data_buf[872] : encrypted_data_buf_next[872];   // modexp_top.v(751)
    assign n8792 = rst ? encrypted_data_buf[871] : encrypted_data_buf_next[871];   // modexp_top.v(751)
    assign n8793 = rst ? encrypted_data_buf[870] : encrypted_data_buf_next[870];   // modexp_top.v(751)
    assign n8794 = rst ? encrypted_data_buf[869] : encrypted_data_buf_next[869];   // modexp_top.v(751)
    assign n8795 = rst ? encrypted_data_buf[868] : encrypted_data_buf_next[868];   // modexp_top.v(751)
    assign n8796 = rst ? encrypted_data_buf[867] : encrypted_data_buf_next[867];   // modexp_top.v(751)
    assign n8797 = rst ? encrypted_data_buf[866] : encrypted_data_buf_next[866];   // modexp_top.v(751)
    assign n8798 = rst ? encrypted_data_buf[865] : encrypted_data_buf_next[865];   // modexp_top.v(751)
    assign n8799 = rst ? encrypted_data_buf[864] : encrypted_data_buf_next[864];   // modexp_top.v(751)
    assign n8800 = rst ? encrypted_data_buf[863] : encrypted_data_buf_next[863];   // modexp_top.v(751)
    assign n8801 = rst ? encrypted_data_buf[862] : encrypted_data_buf_next[862];   // modexp_top.v(751)
    assign n8802 = rst ? encrypted_data_buf[861] : encrypted_data_buf_next[861];   // modexp_top.v(751)
    assign n8803 = rst ? encrypted_data_buf[860] : encrypted_data_buf_next[860];   // modexp_top.v(751)
    assign n8804 = rst ? encrypted_data_buf[859] : encrypted_data_buf_next[859];   // modexp_top.v(751)
    assign n8805 = rst ? encrypted_data_buf[858] : encrypted_data_buf_next[858];   // modexp_top.v(751)
    assign n8806 = rst ? encrypted_data_buf[857] : encrypted_data_buf_next[857];   // modexp_top.v(751)
    assign n8807 = rst ? encrypted_data_buf[856] : encrypted_data_buf_next[856];   // modexp_top.v(751)
    assign n8808 = rst ? encrypted_data_buf[855] : encrypted_data_buf_next[855];   // modexp_top.v(751)
    assign n8809 = rst ? encrypted_data_buf[854] : encrypted_data_buf_next[854];   // modexp_top.v(751)
    assign n8810 = rst ? encrypted_data_buf[853] : encrypted_data_buf_next[853];   // modexp_top.v(751)
    assign n8811 = rst ? encrypted_data_buf[852] : encrypted_data_buf_next[852];   // modexp_top.v(751)
    assign n8812 = rst ? encrypted_data_buf[851] : encrypted_data_buf_next[851];   // modexp_top.v(751)
    assign n8813 = rst ? encrypted_data_buf[850] : encrypted_data_buf_next[850];   // modexp_top.v(751)
    assign n8814 = rst ? encrypted_data_buf[849] : encrypted_data_buf_next[849];   // modexp_top.v(751)
    assign n8815 = rst ? encrypted_data_buf[848] : encrypted_data_buf_next[848];   // modexp_top.v(751)
    assign n8816 = rst ? encrypted_data_buf[847] : encrypted_data_buf_next[847];   // modexp_top.v(751)
    assign n8817 = rst ? encrypted_data_buf[846] : encrypted_data_buf_next[846];   // modexp_top.v(751)
    assign n8818 = rst ? encrypted_data_buf[845] : encrypted_data_buf_next[845];   // modexp_top.v(751)
    assign n8819 = rst ? encrypted_data_buf[844] : encrypted_data_buf_next[844];   // modexp_top.v(751)
    assign n8820 = rst ? encrypted_data_buf[843] : encrypted_data_buf_next[843];   // modexp_top.v(751)
    assign n8821 = rst ? encrypted_data_buf[842] : encrypted_data_buf_next[842];   // modexp_top.v(751)
    assign n8822 = rst ? encrypted_data_buf[841] : encrypted_data_buf_next[841];   // modexp_top.v(751)
    assign n8823 = rst ? encrypted_data_buf[840] : encrypted_data_buf_next[840];   // modexp_top.v(751)
    assign n8824 = rst ? encrypted_data_buf[839] : encrypted_data_buf_next[839];   // modexp_top.v(751)
    assign n8825 = rst ? encrypted_data_buf[838] : encrypted_data_buf_next[838];   // modexp_top.v(751)
    assign n8826 = rst ? encrypted_data_buf[837] : encrypted_data_buf_next[837];   // modexp_top.v(751)
    assign n8827 = rst ? encrypted_data_buf[836] : encrypted_data_buf_next[836];   // modexp_top.v(751)
    assign n8828 = rst ? encrypted_data_buf[835] : encrypted_data_buf_next[835];   // modexp_top.v(751)
    assign n8829 = rst ? encrypted_data_buf[834] : encrypted_data_buf_next[834];   // modexp_top.v(751)
    assign n8830 = rst ? encrypted_data_buf[833] : encrypted_data_buf_next[833];   // modexp_top.v(751)
    assign n8831 = rst ? encrypted_data_buf[832] : encrypted_data_buf_next[832];   // modexp_top.v(751)
    assign n8832 = rst ? encrypted_data_buf[831] : encrypted_data_buf_next[831];   // modexp_top.v(751)
    assign n8833 = rst ? encrypted_data_buf[830] : encrypted_data_buf_next[830];   // modexp_top.v(751)
    assign n8834 = rst ? encrypted_data_buf[829] : encrypted_data_buf_next[829];   // modexp_top.v(751)
    assign n8835 = rst ? encrypted_data_buf[828] : encrypted_data_buf_next[828];   // modexp_top.v(751)
    assign n8836 = rst ? encrypted_data_buf[827] : encrypted_data_buf_next[827];   // modexp_top.v(751)
    assign n8837 = rst ? encrypted_data_buf[826] : encrypted_data_buf_next[826];   // modexp_top.v(751)
    assign n8838 = rst ? encrypted_data_buf[825] : encrypted_data_buf_next[825];   // modexp_top.v(751)
    assign n8839 = rst ? encrypted_data_buf[824] : encrypted_data_buf_next[824];   // modexp_top.v(751)
    assign n8840 = rst ? encrypted_data_buf[823] : encrypted_data_buf_next[823];   // modexp_top.v(751)
    assign n8841 = rst ? encrypted_data_buf[822] : encrypted_data_buf_next[822];   // modexp_top.v(751)
    assign n8842 = rst ? encrypted_data_buf[821] : encrypted_data_buf_next[821];   // modexp_top.v(751)
    assign n8843 = rst ? encrypted_data_buf[820] : encrypted_data_buf_next[820];   // modexp_top.v(751)
    assign n8844 = rst ? encrypted_data_buf[819] : encrypted_data_buf_next[819];   // modexp_top.v(751)
    assign n8845 = rst ? encrypted_data_buf[818] : encrypted_data_buf_next[818];   // modexp_top.v(751)
    assign n8846 = rst ? encrypted_data_buf[817] : encrypted_data_buf_next[817];   // modexp_top.v(751)
    assign n8847 = rst ? encrypted_data_buf[816] : encrypted_data_buf_next[816];   // modexp_top.v(751)
    assign n8848 = rst ? encrypted_data_buf[815] : encrypted_data_buf_next[815];   // modexp_top.v(751)
    assign n8849 = rst ? encrypted_data_buf[814] : encrypted_data_buf_next[814];   // modexp_top.v(751)
    assign n8850 = rst ? encrypted_data_buf[813] : encrypted_data_buf_next[813];   // modexp_top.v(751)
    assign n8851 = rst ? encrypted_data_buf[812] : encrypted_data_buf_next[812];   // modexp_top.v(751)
    assign n8852 = rst ? encrypted_data_buf[811] : encrypted_data_buf_next[811];   // modexp_top.v(751)
    assign n8853 = rst ? encrypted_data_buf[810] : encrypted_data_buf_next[810];   // modexp_top.v(751)
    assign n8854 = rst ? encrypted_data_buf[809] : encrypted_data_buf_next[809];   // modexp_top.v(751)
    assign n8855 = rst ? encrypted_data_buf[808] : encrypted_data_buf_next[808];   // modexp_top.v(751)
    assign n8856 = rst ? encrypted_data_buf[807] : encrypted_data_buf_next[807];   // modexp_top.v(751)
    assign n8857 = rst ? encrypted_data_buf[806] : encrypted_data_buf_next[806];   // modexp_top.v(751)
    assign n8858 = rst ? encrypted_data_buf[805] : encrypted_data_buf_next[805];   // modexp_top.v(751)
    assign n8859 = rst ? encrypted_data_buf[804] : encrypted_data_buf_next[804];   // modexp_top.v(751)
    assign n8860 = rst ? encrypted_data_buf[803] : encrypted_data_buf_next[803];   // modexp_top.v(751)
    assign n8861 = rst ? encrypted_data_buf[802] : encrypted_data_buf_next[802];   // modexp_top.v(751)
    assign n8862 = rst ? encrypted_data_buf[801] : encrypted_data_buf_next[801];   // modexp_top.v(751)
    assign n8863 = rst ? encrypted_data_buf[800] : encrypted_data_buf_next[800];   // modexp_top.v(751)
    assign n8864 = rst ? encrypted_data_buf[799] : encrypted_data_buf_next[799];   // modexp_top.v(751)
    assign n8865 = rst ? encrypted_data_buf[798] : encrypted_data_buf_next[798];   // modexp_top.v(751)
    assign n8866 = rst ? encrypted_data_buf[797] : encrypted_data_buf_next[797];   // modexp_top.v(751)
    assign n8867 = rst ? encrypted_data_buf[796] : encrypted_data_buf_next[796];   // modexp_top.v(751)
    assign n8868 = rst ? encrypted_data_buf[795] : encrypted_data_buf_next[795];   // modexp_top.v(751)
    assign n8869 = rst ? encrypted_data_buf[794] : encrypted_data_buf_next[794];   // modexp_top.v(751)
    assign n8870 = rst ? encrypted_data_buf[793] : encrypted_data_buf_next[793];   // modexp_top.v(751)
    assign n8871 = rst ? encrypted_data_buf[792] : encrypted_data_buf_next[792];   // modexp_top.v(751)
    assign n8872 = rst ? encrypted_data_buf[791] : encrypted_data_buf_next[791];   // modexp_top.v(751)
    assign n8873 = rst ? encrypted_data_buf[790] : encrypted_data_buf_next[790];   // modexp_top.v(751)
    assign n8874 = rst ? encrypted_data_buf[789] : encrypted_data_buf_next[789];   // modexp_top.v(751)
    assign n8875 = rst ? encrypted_data_buf[788] : encrypted_data_buf_next[788];   // modexp_top.v(751)
    assign n8876 = rst ? encrypted_data_buf[787] : encrypted_data_buf_next[787];   // modexp_top.v(751)
    assign n8877 = rst ? encrypted_data_buf[786] : encrypted_data_buf_next[786];   // modexp_top.v(751)
    assign n8878 = rst ? encrypted_data_buf[785] : encrypted_data_buf_next[785];   // modexp_top.v(751)
    assign n8879 = rst ? encrypted_data_buf[784] : encrypted_data_buf_next[784];   // modexp_top.v(751)
    assign n8880 = rst ? encrypted_data_buf[783] : encrypted_data_buf_next[783];   // modexp_top.v(751)
    assign n8881 = rst ? encrypted_data_buf[782] : encrypted_data_buf_next[782];   // modexp_top.v(751)
    assign n8882 = rst ? encrypted_data_buf[781] : encrypted_data_buf_next[781];   // modexp_top.v(751)
    assign n8883 = rst ? encrypted_data_buf[780] : encrypted_data_buf_next[780];   // modexp_top.v(751)
    assign n8884 = rst ? encrypted_data_buf[779] : encrypted_data_buf_next[779];   // modexp_top.v(751)
    assign n8885 = rst ? encrypted_data_buf[778] : encrypted_data_buf_next[778];   // modexp_top.v(751)
    assign n8886 = rst ? encrypted_data_buf[777] : encrypted_data_buf_next[777];   // modexp_top.v(751)
    assign n8887 = rst ? encrypted_data_buf[776] : encrypted_data_buf_next[776];   // modexp_top.v(751)
    assign n8888 = rst ? encrypted_data_buf[775] : encrypted_data_buf_next[775];   // modexp_top.v(751)
    assign n8889 = rst ? encrypted_data_buf[774] : encrypted_data_buf_next[774];   // modexp_top.v(751)
    assign n8890 = rst ? encrypted_data_buf[773] : encrypted_data_buf_next[773];   // modexp_top.v(751)
    assign n8891 = rst ? encrypted_data_buf[772] : encrypted_data_buf_next[772];   // modexp_top.v(751)
    assign n8892 = rst ? encrypted_data_buf[771] : encrypted_data_buf_next[771];   // modexp_top.v(751)
    assign n8893 = rst ? encrypted_data_buf[770] : encrypted_data_buf_next[770];   // modexp_top.v(751)
    assign n8894 = rst ? encrypted_data_buf[769] : encrypted_data_buf_next[769];   // modexp_top.v(751)
    assign n8895 = rst ? encrypted_data_buf[768] : encrypted_data_buf_next[768];   // modexp_top.v(751)
    assign n8896 = rst ? encrypted_data_buf[767] : encrypted_data_buf_next[767];   // modexp_top.v(751)
    assign n8897 = rst ? encrypted_data_buf[766] : encrypted_data_buf_next[766];   // modexp_top.v(751)
    assign n8898 = rst ? encrypted_data_buf[765] : encrypted_data_buf_next[765];   // modexp_top.v(751)
    assign n8899 = rst ? encrypted_data_buf[764] : encrypted_data_buf_next[764];   // modexp_top.v(751)
    assign n8900 = rst ? encrypted_data_buf[763] : encrypted_data_buf_next[763];   // modexp_top.v(751)
    assign n8901 = rst ? encrypted_data_buf[762] : encrypted_data_buf_next[762];   // modexp_top.v(751)
    assign n8902 = rst ? encrypted_data_buf[761] : encrypted_data_buf_next[761];   // modexp_top.v(751)
    assign n8903 = rst ? encrypted_data_buf[760] : encrypted_data_buf_next[760];   // modexp_top.v(751)
    assign n8904 = rst ? encrypted_data_buf[759] : encrypted_data_buf_next[759];   // modexp_top.v(751)
    assign n8905 = rst ? encrypted_data_buf[758] : encrypted_data_buf_next[758];   // modexp_top.v(751)
    assign n8906 = rst ? encrypted_data_buf[757] : encrypted_data_buf_next[757];   // modexp_top.v(751)
    assign n8907 = rst ? encrypted_data_buf[756] : encrypted_data_buf_next[756];   // modexp_top.v(751)
    assign n8908 = rst ? encrypted_data_buf[755] : encrypted_data_buf_next[755];   // modexp_top.v(751)
    assign n8909 = rst ? encrypted_data_buf[754] : encrypted_data_buf_next[754];   // modexp_top.v(751)
    assign n8910 = rst ? encrypted_data_buf[753] : encrypted_data_buf_next[753];   // modexp_top.v(751)
    assign n8911 = rst ? encrypted_data_buf[752] : encrypted_data_buf_next[752];   // modexp_top.v(751)
    assign n8912 = rst ? encrypted_data_buf[751] : encrypted_data_buf_next[751];   // modexp_top.v(751)
    assign n8913 = rst ? encrypted_data_buf[750] : encrypted_data_buf_next[750];   // modexp_top.v(751)
    assign n8914 = rst ? encrypted_data_buf[749] : encrypted_data_buf_next[749];   // modexp_top.v(751)
    assign n8915 = rst ? encrypted_data_buf[748] : encrypted_data_buf_next[748];   // modexp_top.v(751)
    assign n8916 = rst ? encrypted_data_buf[747] : encrypted_data_buf_next[747];   // modexp_top.v(751)
    assign n8917 = rst ? encrypted_data_buf[746] : encrypted_data_buf_next[746];   // modexp_top.v(751)
    assign n8918 = rst ? encrypted_data_buf[745] : encrypted_data_buf_next[745];   // modexp_top.v(751)
    assign n8919 = rst ? encrypted_data_buf[744] : encrypted_data_buf_next[744];   // modexp_top.v(751)
    assign n8920 = rst ? encrypted_data_buf[743] : encrypted_data_buf_next[743];   // modexp_top.v(751)
    assign n8921 = rst ? encrypted_data_buf[742] : encrypted_data_buf_next[742];   // modexp_top.v(751)
    assign n8922 = rst ? encrypted_data_buf[741] : encrypted_data_buf_next[741];   // modexp_top.v(751)
    assign n8923 = rst ? encrypted_data_buf[740] : encrypted_data_buf_next[740];   // modexp_top.v(751)
    assign n8924 = rst ? encrypted_data_buf[739] : encrypted_data_buf_next[739];   // modexp_top.v(751)
    assign n8925 = rst ? encrypted_data_buf[738] : encrypted_data_buf_next[738];   // modexp_top.v(751)
    assign n8926 = rst ? encrypted_data_buf[737] : encrypted_data_buf_next[737];   // modexp_top.v(751)
    assign n8927 = rst ? encrypted_data_buf[736] : encrypted_data_buf_next[736];   // modexp_top.v(751)
    assign n8928 = rst ? encrypted_data_buf[735] : encrypted_data_buf_next[735];   // modexp_top.v(751)
    assign n8929 = rst ? encrypted_data_buf[734] : encrypted_data_buf_next[734];   // modexp_top.v(751)
    assign n8930 = rst ? encrypted_data_buf[733] : encrypted_data_buf_next[733];   // modexp_top.v(751)
    assign n8931 = rst ? encrypted_data_buf[732] : encrypted_data_buf_next[732];   // modexp_top.v(751)
    assign n8932 = rst ? encrypted_data_buf[731] : encrypted_data_buf_next[731];   // modexp_top.v(751)
    assign n8933 = rst ? encrypted_data_buf[730] : encrypted_data_buf_next[730];   // modexp_top.v(751)
    assign n8934 = rst ? encrypted_data_buf[729] : encrypted_data_buf_next[729];   // modexp_top.v(751)
    assign n8935 = rst ? encrypted_data_buf[728] : encrypted_data_buf_next[728];   // modexp_top.v(751)
    assign n8936 = rst ? encrypted_data_buf[727] : encrypted_data_buf_next[727];   // modexp_top.v(751)
    assign n8937 = rst ? encrypted_data_buf[726] : encrypted_data_buf_next[726];   // modexp_top.v(751)
    assign n8938 = rst ? encrypted_data_buf[725] : encrypted_data_buf_next[725];   // modexp_top.v(751)
    assign n8939 = rst ? encrypted_data_buf[724] : encrypted_data_buf_next[724];   // modexp_top.v(751)
    assign n8940 = rst ? encrypted_data_buf[723] : encrypted_data_buf_next[723];   // modexp_top.v(751)
    assign n8941 = rst ? encrypted_data_buf[722] : encrypted_data_buf_next[722];   // modexp_top.v(751)
    assign n8942 = rst ? encrypted_data_buf[721] : encrypted_data_buf_next[721];   // modexp_top.v(751)
    assign n8943 = rst ? encrypted_data_buf[720] : encrypted_data_buf_next[720];   // modexp_top.v(751)
    assign n8944 = rst ? encrypted_data_buf[719] : encrypted_data_buf_next[719];   // modexp_top.v(751)
    assign n8945 = rst ? encrypted_data_buf[718] : encrypted_data_buf_next[718];   // modexp_top.v(751)
    assign n8946 = rst ? encrypted_data_buf[717] : encrypted_data_buf_next[717];   // modexp_top.v(751)
    assign n8947 = rst ? encrypted_data_buf[716] : encrypted_data_buf_next[716];   // modexp_top.v(751)
    assign n8948 = rst ? encrypted_data_buf[715] : encrypted_data_buf_next[715];   // modexp_top.v(751)
    assign n8949 = rst ? encrypted_data_buf[714] : encrypted_data_buf_next[714];   // modexp_top.v(751)
    assign n8950 = rst ? encrypted_data_buf[713] : encrypted_data_buf_next[713];   // modexp_top.v(751)
    assign n8951 = rst ? encrypted_data_buf[712] : encrypted_data_buf_next[712];   // modexp_top.v(751)
    assign n8952 = rst ? encrypted_data_buf[711] : encrypted_data_buf_next[711];   // modexp_top.v(751)
    assign n8953 = rst ? encrypted_data_buf[710] : encrypted_data_buf_next[710];   // modexp_top.v(751)
    assign n8954 = rst ? encrypted_data_buf[709] : encrypted_data_buf_next[709];   // modexp_top.v(751)
    assign n8955 = rst ? encrypted_data_buf[708] : encrypted_data_buf_next[708];   // modexp_top.v(751)
    assign n8956 = rst ? encrypted_data_buf[707] : encrypted_data_buf_next[707];   // modexp_top.v(751)
    assign n8957 = rst ? encrypted_data_buf[706] : encrypted_data_buf_next[706];   // modexp_top.v(751)
    assign n8958 = rst ? encrypted_data_buf[705] : encrypted_data_buf_next[705];   // modexp_top.v(751)
    assign n8959 = rst ? encrypted_data_buf[704] : encrypted_data_buf_next[704];   // modexp_top.v(751)
    assign n8960 = rst ? encrypted_data_buf[703] : encrypted_data_buf_next[703];   // modexp_top.v(751)
    assign n8961 = rst ? encrypted_data_buf[702] : encrypted_data_buf_next[702];   // modexp_top.v(751)
    assign n8962 = rst ? encrypted_data_buf[701] : encrypted_data_buf_next[701];   // modexp_top.v(751)
    assign n8963 = rst ? encrypted_data_buf[700] : encrypted_data_buf_next[700];   // modexp_top.v(751)
    assign n8964 = rst ? encrypted_data_buf[699] : encrypted_data_buf_next[699];   // modexp_top.v(751)
    assign n8965 = rst ? encrypted_data_buf[698] : encrypted_data_buf_next[698];   // modexp_top.v(751)
    assign n8966 = rst ? encrypted_data_buf[697] : encrypted_data_buf_next[697];   // modexp_top.v(751)
    assign n8967 = rst ? encrypted_data_buf[696] : encrypted_data_buf_next[696];   // modexp_top.v(751)
    assign n8968 = rst ? encrypted_data_buf[695] : encrypted_data_buf_next[695];   // modexp_top.v(751)
    assign n8969 = rst ? encrypted_data_buf[694] : encrypted_data_buf_next[694];   // modexp_top.v(751)
    assign n8970 = rst ? encrypted_data_buf[693] : encrypted_data_buf_next[693];   // modexp_top.v(751)
    assign n8971 = rst ? encrypted_data_buf[692] : encrypted_data_buf_next[692];   // modexp_top.v(751)
    assign n8972 = rst ? encrypted_data_buf[691] : encrypted_data_buf_next[691];   // modexp_top.v(751)
    assign n8973 = rst ? encrypted_data_buf[690] : encrypted_data_buf_next[690];   // modexp_top.v(751)
    assign n8974 = rst ? encrypted_data_buf[689] : encrypted_data_buf_next[689];   // modexp_top.v(751)
    assign n8975 = rst ? encrypted_data_buf[688] : encrypted_data_buf_next[688];   // modexp_top.v(751)
    assign n8976 = rst ? encrypted_data_buf[687] : encrypted_data_buf_next[687];   // modexp_top.v(751)
    assign n8977 = rst ? encrypted_data_buf[686] : encrypted_data_buf_next[686];   // modexp_top.v(751)
    assign n8978 = rst ? encrypted_data_buf[685] : encrypted_data_buf_next[685];   // modexp_top.v(751)
    assign n8979 = rst ? encrypted_data_buf[684] : encrypted_data_buf_next[684];   // modexp_top.v(751)
    assign n8980 = rst ? encrypted_data_buf[683] : encrypted_data_buf_next[683];   // modexp_top.v(751)
    assign n8981 = rst ? encrypted_data_buf[682] : encrypted_data_buf_next[682];   // modexp_top.v(751)
    assign n8982 = rst ? encrypted_data_buf[681] : encrypted_data_buf_next[681];   // modexp_top.v(751)
    assign n8983 = rst ? encrypted_data_buf[680] : encrypted_data_buf_next[680];   // modexp_top.v(751)
    assign n8984 = rst ? encrypted_data_buf[679] : encrypted_data_buf_next[679];   // modexp_top.v(751)
    assign n8985 = rst ? encrypted_data_buf[678] : encrypted_data_buf_next[678];   // modexp_top.v(751)
    assign n8986 = rst ? encrypted_data_buf[677] : encrypted_data_buf_next[677];   // modexp_top.v(751)
    assign n8987 = rst ? encrypted_data_buf[676] : encrypted_data_buf_next[676];   // modexp_top.v(751)
    assign n8988 = rst ? encrypted_data_buf[675] : encrypted_data_buf_next[675];   // modexp_top.v(751)
    assign n8989 = rst ? encrypted_data_buf[674] : encrypted_data_buf_next[674];   // modexp_top.v(751)
    assign n8990 = rst ? encrypted_data_buf[673] : encrypted_data_buf_next[673];   // modexp_top.v(751)
    assign n8991 = rst ? encrypted_data_buf[672] : encrypted_data_buf_next[672];   // modexp_top.v(751)
    assign n8992 = rst ? encrypted_data_buf[671] : encrypted_data_buf_next[671];   // modexp_top.v(751)
    assign n8993 = rst ? encrypted_data_buf[670] : encrypted_data_buf_next[670];   // modexp_top.v(751)
    assign n8994 = rst ? encrypted_data_buf[669] : encrypted_data_buf_next[669];   // modexp_top.v(751)
    assign n8995 = rst ? encrypted_data_buf[668] : encrypted_data_buf_next[668];   // modexp_top.v(751)
    assign n8996 = rst ? encrypted_data_buf[667] : encrypted_data_buf_next[667];   // modexp_top.v(751)
    assign n8997 = rst ? encrypted_data_buf[666] : encrypted_data_buf_next[666];   // modexp_top.v(751)
    assign n8998 = rst ? encrypted_data_buf[665] : encrypted_data_buf_next[665];   // modexp_top.v(751)
    assign n8999 = rst ? encrypted_data_buf[664] : encrypted_data_buf_next[664];   // modexp_top.v(751)
    assign n9000 = rst ? encrypted_data_buf[663] : encrypted_data_buf_next[663];   // modexp_top.v(751)
    assign n9001 = rst ? encrypted_data_buf[662] : encrypted_data_buf_next[662];   // modexp_top.v(751)
    assign n9002 = rst ? encrypted_data_buf[661] : encrypted_data_buf_next[661];   // modexp_top.v(751)
    assign n9003 = rst ? encrypted_data_buf[660] : encrypted_data_buf_next[660];   // modexp_top.v(751)
    assign n9004 = rst ? encrypted_data_buf[659] : encrypted_data_buf_next[659];   // modexp_top.v(751)
    assign n9005 = rst ? encrypted_data_buf[658] : encrypted_data_buf_next[658];   // modexp_top.v(751)
    assign n9006 = rst ? encrypted_data_buf[657] : encrypted_data_buf_next[657];   // modexp_top.v(751)
    assign n9007 = rst ? encrypted_data_buf[656] : encrypted_data_buf_next[656];   // modexp_top.v(751)
    assign n9008 = rst ? encrypted_data_buf[655] : encrypted_data_buf_next[655];   // modexp_top.v(751)
    assign n9009 = rst ? encrypted_data_buf[654] : encrypted_data_buf_next[654];   // modexp_top.v(751)
    assign n9010 = rst ? encrypted_data_buf[653] : encrypted_data_buf_next[653];   // modexp_top.v(751)
    assign n9011 = rst ? encrypted_data_buf[652] : encrypted_data_buf_next[652];   // modexp_top.v(751)
    assign n9012 = rst ? encrypted_data_buf[651] : encrypted_data_buf_next[651];   // modexp_top.v(751)
    assign n9013 = rst ? encrypted_data_buf[650] : encrypted_data_buf_next[650];   // modexp_top.v(751)
    assign n9014 = rst ? encrypted_data_buf[649] : encrypted_data_buf_next[649];   // modexp_top.v(751)
    assign n9015 = rst ? encrypted_data_buf[648] : encrypted_data_buf_next[648];   // modexp_top.v(751)
    assign n9016 = rst ? encrypted_data_buf[647] : encrypted_data_buf_next[647];   // modexp_top.v(751)
    assign n9017 = rst ? encrypted_data_buf[646] : encrypted_data_buf_next[646];   // modexp_top.v(751)
    assign n9018 = rst ? encrypted_data_buf[645] : encrypted_data_buf_next[645];   // modexp_top.v(751)
    assign n9019 = rst ? encrypted_data_buf[644] : encrypted_data_buf_next[644];   // modexp_top.v(751)
    assign n9020 = rst ? encrypted_data_buf[643] : encrypted_data_buf_next[643];   // modexp_top.v(751)
    assign n9021 = rst ? encrypted_data_buf[642] : encrypted_data_buf_next[642];   // modexp_top.v(751)
    assign n9022 = rst ? encrypted_data_buf[641] : encrypted_data_buf_next[641];   // modexp_top.v(751)
    assign n9023 = rst ? encrypted_data_buf[640] : encrypted_data_buf_next[640];   // modexp_top.v(751)
    assign n9024 = rst ? encrypted_data_buf[639] : encrypted_data_buf_next[639];   // modexp_top.v(751)
    assign n9025 = rst ? encrypted_data_buf[638] : encrypted_data_buf_next[638];   // modexp_top.v(751)
    assign n9026 = rst ? encrypted_data_buf[637] : encrypted_data_buf_next[637];   // modexp_top.v(751)
    assign n9027 = rst ? encrypted_data_buf[636] : encrypted_data_buf_next[636];   // modexp_top.v(751)
    assign n9028 = rst ? encrypted_data_buf[635] : encrypted_data_buf_next[635];   // modexp_top.v(751)
    assign n9029 = rst ? encrypted_data_buf[634] : encrypted_data_buf_next[634];   // modexp_top.v(751)
    assign n9030 = rst ? encrypted_data_buf[633] : encrypted_data_buf_next[633];   // modexp_top.v(751)
    assign n9031 = rst ? encrypted_data_buf[632] : encrypted_data_buf_next[632];   // modexp_top.v(751)
    assign n9032 = rst ? encrypted_data_buf[631] : encrypted_data_buf_next[631];   // modexp_top.v(751)
    assign n9033 = rst ? encrypted_data_buf[630] : encrypted_data_buf_next[630];   // modexp_top.v(751)
    assign n9034 = rst ? encrypted_data_buf[629] : encrypted_data_buf_next[629];   // modexp_top.v(751)
    assign n9035 = rst ? encrypted_data_buf[628] : encrypted_data_buf_next[628];   // modexp_top.v(751)
    assign n9036 = rst ? encrypted_data_buf[627] : encrypted_data_buf_next[627];   // modexp_top.v(751)
    assign n9037 = rst ? encrypted_data_buf[626] : encrypted_data_buf_next[626];   // modexp_top.v(751)
    assign n9038 = rst ? encrypted_data_buf[625] : encrypted_data_buf_next[625];   // modexp_top.v(751)
    assign n9039 = rst ? encrypted_data_buf[624] : encrypted_data_buf_next[624];   // modexp_top.v(751)
    assign n9040 = rst ? encrypted_data_buf[623] : encrypted_data_buf_next[623];   // modexp_top.v(751)
    assign n9041 = rst ? encrypted_data_buf[622] : encrypted_data_buf_next[622];   // modexp_top.v(751)
    assign n9042 = rst ? encrypted_data_buf[621] : encrypted_data_buf_next[621];   // modexp_top.v(751)
    assign n9043 = rst ? encrypted_data_buf[620] : encrypted_data_buf_next[620];   // modexp_top.v(751)
    assign n9044 = rst ? encrypted_data_buf[619] : encrypted_data_buf_next[619];   // modexp_top.v(751)
    assign n9045 = rst ? encrypted_data_buf[618] : encrypted_data_buf_next[618];   // modexp_top.v(751)
    assign n9046 = rst ? encrypted_data_buf[617] : encrypted_data_buf_next[617];   // modexp_top.v(751)
    assign n9047 = rst ? encrypted_data_buf[616] : encrypted_data_buf_next[616];   // modexp_top.v(751)
    assign n9048 = rst ? encrypted_data_buf[615] : encrypted_data_buf_next[615];   // modexp_top.v(751)
    assign n9049 = rst ? encrypted_data_buf[614] : encrypted_data_buf_next[614];   // modexp_top.v(751)
    assign n9050 = rst ? encrypted_data_buf[613] : encrypted_data_buf_next[613];   // modexp_top.v(751)
    assign n9051 = rst ? encrypted_data_buf[612] : encrypted_data_buf_next[612];   // modexp_top.v(751)
    assign n9052 = rst ? encrypted_data_buf[611] : encrypted_data_buf_next[611];   // modexp_top.v(751)
    assign n9053 = rst ? encrypted_data_buf[610] : encrypted_data_buf_next[610];   // modexp_top.v(751)
    assign n9054 = rst ? encrypted_data_buf[609] : encrypted_data_buf_next[609];   // modexp_top.v(751)
    assign n9055 = rst ? encrypted_data_buf[608] : encrypted_data_buf_next[608];   // modexp_top.v(751)
    assign n9056 = rst ? encrypted_data_buf[607] : encrypted_data_buf_next[607];   // modexp_top.v(751)
    assign n9057 = rst ? encrypted_data_buf[606] : encrypted_data_buf_next[606];   // modexp_top.v(751)
    assign n9058 = rst ? encrypted_data_buf[605] : encrypted_data_buf_next[605];   // modexp_top.v(751)
    assign n9059 = rst ? encrypted_data_buf[604] : encrypted_data_buf_next[604];   // modexp_top.v(751)
    assign n9060 = rst ? encrypted_data_buf[603] : encrypted_data_buf_next[603];   // modexp_top.v(751)
    assign n9061 = rst ? encrypted_data_buf[602] : encrypted_data_buf_next[602];   // modexp_top.v(751)
    assign n9062 = rst ? encrypted_data_buf[601] : encrypted_data_buf_next[601];   // modexp_top.v(751)
    assign n9063 = rst ? encrypted_data_buf[600] : encrypted_data_buf_next[600];   // modexp_top.v(751)
    assign n9064 = rst ? encrypted_data_buf[599] : encrypted_data_buf_next[599];   // modexp_top.v(751)
    assign n9065 = rst ? encrypted_data_buf[598] : encrypted_data_buf_next[598];   // modexp_top.v(751)
    assign n9066 = rst ? encrypted_data_buf[597] : encrypted_data_buf_next[597];   // modexp_top.v(751)
    assign n9067 = rst ? encrypted_data_buf[596] : encrypted_data_buf_next[596];   // modexp_top.v(751)
    assign n9068 = rst ? encrypted_data_buf[595] : encrypted_data_buf_next[595];   // modexp_top.v(751)
    assign n9069 = rst ? encrypted_data_buf[594] : encrypted_data_buf_next[594];   // modexp_top.v(751)
    assign n9070 = rst ? encrypted_data_buf[593] : encrypted_data_buf_next[593];   // modexp_top.v(751)
    assign n9071 = rst ? encrypted_data_buf[592] : encrypted_data_buf_next[592];   // modexp_top.v(751)
    assign n9072 = rst ? encrypted_data_buf[591] : encrypted_data_buf_next[591];   // modexp_top.v(751)
    assign n9073 = rst ? encrypted_data_buf[590] : encrypted_data_buf_next[590];   // modexp_top.v(751)
    assign n9074 = rst ? encrypted_data_buf[589] : encrypted_data_buf_next[589];   // modexp_top.v(751)
    assign n9075 = rst ? encrypted_data_buf[588] : encrypted_data_buf_next[588];   // modexp_top.v(751)
    assign n9076 = rst ? encrypted_data_buf[587] : encrypted_data_buf_next[587];   // modexp_top.v(751)
    assign n9077 = rst ? encrypted_data_buf[586] : encrypted_data_buf_next[586];   // modexp_top.v(751)
    assign n9078 = rst ? encrypted_data_buf[585] : encrypted_data_buf_next[585];   // modexp_top.v(751)
    assign n9079 = rst ? encrypted_data_buf[584] : encrypted_data_buf_next[584];   // modexp_top.v(751)
    assign n9080 = rst ? encrypted_data_buf[583] : encrypted_data_buf_next[583];   // modexp_top.v(751)
    assign n9081 = rst ? encrypted_data_buf[582] : encrypted_data_buf_next[582];   // modexp_top.v(751)
    assign n9082 = rst ? encrypted_data_buf[581] : encrypted_data_buf_next[581];   // modexp_top.v(751)
    assign n9083 = rst ? encrypted_data_buf[580] : encrypted_data_buf_next[580];   // modexp_top.v(751)
    assign n9084 = rst ? encrypted_data_buf[579] : encrypted_data_buf_next[579];   // modexp_top.v(751)
    assign n9085 = rst ? encrypted_data_buf[578] : encrypted_data_buf_next[578];   // modexp_top.v(751)
    assign n9086 = rst ? encrypted_data_buf[577] : encrypted_data_buf_next[577];   // modexp_top.v(751)
    assign n9087 = rst ? encrypted_data_buf[576] : encrypted_data_buf_next[576];   // modexp_top.v(751)
    assign n9088 = rst ? encrypted_data_buf[575] : encrypted_data_buf_next[575];   // modexp_top.v(751)
    assign n9089 = rst ? encrypted_data_buf[574] : encrypted_data_buf_next[574];   // modexp_top.v(751)
    assign n9090 = rst ? encrypted_data_buf[573] : encrypted_data_buf_next[573];   // modexp_top.v(751)
    assign n9091 = rst ? encrypted_data_buf[572] : encrypted_data_buf_next[572];   // modexp_top.v(751)
    assign n9092 = rst ? encrypted_data_buf[571] : encrypted_data_buf_next[571];   // modexp_top.v(751)
    assign n9093 = rst ? encrypted_data_buf[570] : encrypted_data_buf_next[570];   // modexp_top.v(751)
    assign n9094 = rst ? encrypted_data_buf[569] : encrypted_data_buf_next[569];   // modexp_top.v(751)
    assign n9095 = rst ? encrypted_data_buf[568] : encrypted_data_buf_next[568];   // modexp_top.v(751)
    assign n9096 = rst ? encrypted_data_buf[567] : encrypted_data_buf_next[567];   // modexp_top.v(751)
    assign n9097 = rst ? encrypted_data_buf[566] : encrypted_data_buf_next[566];   // modexp_top.v(751)
    assign n9098 = rst ? encrypted_data_buf[565] : encrypted_data_buf_next[565];   // modexp_top.v(751)
    assign n9099 = rst ? encrypted_data_buf[564] : encrypted_data_buf_next[564];   // modexp_top.v(751)
    assign n9100 = rst ? encrypted_data_buf[563] : encrypted_data_buf_next[563];   // modexp_top.v(751)
    assign n9101 = rst ? encrypted_data_buf[562] : encrypted_data_buf_next[562];   // modexp_top.v(751)
    assign n9102 = rst ? encrypted_data_buf[561] : encrypted_data_buf_next[561];   // modexp_top.v(751)
    assign n9103 = rst ? encrypted_data_buf[560] : encrypted_data_buf_next[560];   // modexp_top.v(751)
    assign n9104 = rst ? encrypted_data_buf[559] : encrypted_data_buf_next[559];   // modexp_top.v(751)
    assign n9105 = rst ? encrypted_data_buf[558] : encrypted_data_buf_next[558];   // modexp_top.v(751)
    assign n9106 = rst ? encrypted_data_buf[557] : encrypted_data_buf_next[557];   // modexp_top.v(751)
    assign n9107 = rst ? encrypted_data_buf[556] : encrypted_data_buf_next[556];   // modexp_top.v(751)
    assign n9108 = rst ? encrypted_data_buf[555] : encrypted_data_buf_next[555];   // modexp_top.v(751)
    assign n9109 = rst ? encrypted_data_buf[554] : encrypted_data_buf_next[554];   // modexp_top.v(751)
    assign n9110 = rst ? encrypted_data_buf[553] : encrypted_data_buf_next[553];   // modexp_top.v(751)
    assign n9111 = rst ? encrypted_data_buf[552] : encrypted_data_buf_next[552];   // modexp_top.v(751)
    assign n9112 = rst ? encrypted_data_buf[551] : encrypted_data_buf_next[551];   // modexp_top.v(751)
    assign n9113 = rst ? encrypted_data_buf[550] : encrypted_data_buf_next[550];   // modexp_top.v(751)
    assign n9114 = rst ? encrypted_data_buf[549] : encrypted_data_buf_next[549];   // modexp_top.v(751)
    assign n9115 = rst ? encrypted_data_buf[548] : encrypted_data_buf_next[548];   // modexp_top.v(751)
    assign n9116 = rst ? encrypted_data_buf[547] : encrypted_data_buf_next[547];   // modexp_top.v(751)
    assign n9117 = rst ? encrypted_data_buf[546] : encrypted_data_buf_next[546];   // modexp_top.v(751)
    assign n9118 = rst ? encrypted_data_buf[545] : encrypted_data_buf_next[545];   // modexp_top.v(751)
    assign n9119 = rst ? encrypted_data_buf[544] : encrypted_data_buf_next[544];   // modexp_top.v(751)
    assign n9120 = rst ? encrypted_data_buf[543] : encrypted_data_buf_next[543];   // modexp_top.v(751)
    assign n9121 = rst ? encrypted_data_buf[542] : encrypted_data_buf_next[542];   // modexp_top.v(751)
    assign n9122 = rst ? encrypted_data_buf[541] : encrypted_data_buf_next[541];   // modexp_top.v(751)
    assign n9123 = rst ? encrypted_data_buf[540] : encrypted_data_buf_next[540];   // modexp_top.v(751)
    assign n9124 = rst ? encrypted_data_buf[539] : encrypted_data_buf_next[539];   // modexp_top.v(751)
    assign n9125 = rst ? encrypted_data_buf[538] : encrypted_data_buf_next[538];   // modexp_top.v(751)
    assign n9126 = rst ? encrypted_data_buf[537] : encrypted_data_buf_next[537];   // modexp_top.v(751)
    assign n9127 = rst ? encrypted_data_buf[536] : encrypted_data_buf_next[536];   // modexp_top.v(751)
    assign n9128 = rst ? encrypted_data_buf[535] : encrypted_data_buf_next[535];   // modexp_top.v(751)
    assign n9129 = rst ? encrypted_data_buf[534] : encrypted_data_buf_next[534];   // modexp_top.v(751)
    assign n9130 = rst ? encrypted_data_buf[533] : encrypted_data_buf_next[533];   // modexp_top.v(751)
    assign n9131 = rst ? encrypted_data_buf[532] : encrypted_data_buf_next[532];   // modexp_top.v(751)
    assign n9132 = rst ? encrypted_data_buf[531] : encrypted_data_buf_next[531];   // modexp_top.v(751)
    assign n9133 = rst ? encrypted_data_buf[530] : encrypted_data_buf_next[530];   // modexp_top.v(751)
    assign n9134 = rst ? encrypted_data_buf[529] : encrypted_data_buf_next[529];   // modexp_top.v(751)
    assign n9135 = rst ? encrypted_data_buf[528] : encrypted_data_buf_next[528];   // modexp_top.v(751)
    assign n9136 = rst ? encrypted_data_buf[527] : encrypted_data_buf_next[527];   // modexp_top.v(751)
    assign n9137 = rst ? encrypted_data_buf[526] : encrypted_data_buf_next[526];   // modexp_top.v(751)
    assign n9138 = rst ? encrypted_data_buf[525] : encrypted_data_buf_next[525];   // modexp_top.v(751)
    assign n9139 = rst ? encrypted_data_buf[524] : encrypted_data_buf_next[524];   // modexp_top.v(751)
    assign n9140 = rst ? encrypted_data_buf[523] : encrypted_data_buf_next[523];   // modexp_top.v(751)
    assign n9141 = rst ? encrypted_data_buf[522] : encrypted_data_buf_next[522];   // modexp_top.v(751)
    assign n9142 = rst ? encrypted_data_buf[521] : encrypted_data_buf_next[521];   // modexp_top.v(751)
    assign n9143 = rst ? encrypted_data_buf[520] : encrypted_data_buf_next[520];   // modexp_top.v(751)
    assign n9144 = rst ? encrypted_data_buf[519] : encrypted_data_buf_next[519];   // modexp_top.v(751)
    assign n9145 = rst ? encrypted_data_buf[518] : encrypted_data_buf_next[518];   // modexp_top.v(751)
    assign n9146 = rst ? encrypted_data_buf[517] : encrypted_data_buf_next[517];   // modexp_top.v(751)
    assign n9147 = rst ? encrypted_data_buf[516] : encrypted_data_buf_next[516];   // modexp_top.v(751)
    assign n9148 = rst ? encrypted_data_buf[515] : encrypted_data_buf_next[515];   // modexp_top.v(751)
    assign n9149 = rst ? encrypted_data_buf[514] : encrypted_data_buf_next[514];   // modexp_top.v(751)
    assign n9150 = rst ? encrypted_data_buf[513] : encrypted_data_buf_next[513];   // modexp_top.v(751)
    assign n9151 = rst ? encrypted_data_buf[512] : encrypted_data_buf_next[512];   // modexp_top.v(751)
    assign n9152 = rst ? encrypted_data_buf[511] : encrypted_data_buf_next[511];   // modexp_top.v(751)
    assign n9153 = rst ? encrypted_data_buf[510] : encrypted_data_buf_next[510];   // modexp_top.v(751)
    assign n9154 = rst ? encrypted_data_buf[509] : encrypted_data_buf_next[509];   // modexp_top.v(751)
    assign n9155 = rst ? encrypted_data_buf[508] : encrypted_data_buf_next[508];   // modexp_top.v(751)
    assign n9156 = rst ? encrypted_data_buf[507] : encrypted_data_buf_next[507];   // modexp_top.v(751)
    assign n9157 = rst ? encrypted_data_buf[506] : encrypted_data_buf_next[506];   // modexp_top.v(751)
    assign n9158 = rst ? encrypted_data_buf[505] : encrypted_data_buf_next[505];   // modexp_top.v(751)
    assign n9159 = rst ? encrypted_data_buf[504] : encrypted_data_buf_next[504];   // modexp_top.v(751)
    assign n9160 = rst ? encrypted_data_buf[503] : encrypted_data_buf_next[503];   // modexp_top.v(751)
    assign n9161 = rst ? encrypted_data_buf[502] : encrypted_data_buf_next[502];   // modexp_top.v(751)
    assign n9162 = rst ? encrypted_data_buf[501] : encrypted_data_buf_next[501];   // modexp_top.v(751)
    assign n9163 = rst ? encrypted_data_buf[500] : encrypted_data_buf_next[500];   // modexp_top.v(751)
    assign n9164 = rst ? encrypted_data_buf[499] : encrypted_data_buf_next[499];   // modexp_top.v(751)
    assign n9165 = rst ? encrypted_data_buf[498] : encrypted_data_buf_next[498];   // modexp_top.v(751)
    assign n9166 = rst ? encrypted_data_buf[497] : encrypted_data_buf_next[497];   // modexp_top.v(751)
    assign n9167 = rst ? encrypted_data_buf[496] : encrypted_data_buf_next[496];   // modexp_top.v(751)
    assign n9168 = rst ? encrypted_data_buf[495] : encrypted_data_buf_next[495];   // modexp_top.v(751)
    assign n9169 = rst ? encrypted_data_buf[494] : encrypted_data_buf_next[494];   // modexp_top.v(751)
    assign n9170 = rst ? encrypted_data_buf[493] : encrypted_data_buf_next[493];   // modexp_top.v(751)
    assign n9171 = rst ? encrypted_data_buf[492] : encrypted_data_buf_next[492];   // modexp_top.v(751)
    assign n9172 = rst ? encrypted_data_buf[491] : encrypted_data_buf_next[491];   // modexp_top.v(751)
    assign n9173 = rst ? encrypted_data_buf[490] : encrypted_data_buf_next[490];   // modexp_top.v(751)
    assign n9174 = rst ? encrypted_data_buf[489] : encrypted_data_buf_next[489];   // modexp_top.v(751)
    assign n9175 = rst ? encrypted_data_buf[488] : encrypted_data_buf_next[488];   // modexp_top.v(751)
    assign n9176 = rst ? encrypted_data_buf[487] : encrypted_data_buf_next[487];   // modexp_top.v(751)
    assign n9177 = rst ? encrypted_data_buf[486] : encrypted_data_buf_next[486];   // modexp_top.v(751)
    assign n9178 = rst ? encrypted_data_buf[485] : encrypted_data_buf_next[485];   // modexp_top.v(751)
    assign n9179 = rst ? encrypted_data_buf[484] : encrypted_data_buf_next[484];   // modexp_top.v(751)
    assign n9180 = rst ? encrypted_data_buf[483] : encrypted_data_buf_next[483];   // modexp_top.v(751)
    assign n9181 = rst ? encrypted_data_buf[482] : encrypted_data_buf_next[482];   // modexp_top.v(751)
    assign n9182 = rst ? encrypted_data_buf[481] : encrypted_data_buf_next[481];   // modexp_top.v(751)
    assign n9183 = rst ? encrypted_data_buf[480] : encrypted_data_buf_next[480];   // modexp_top.v(751)
    assign n9184 = rst ? encrypted_data_buf[479] : encrypted_data_buf_next[479];   // modexp_top.v(751)
    assign n9185 = rst ? encrypted_data_buf[478] : encrypted_data_buf_next[478];   // modexp_top.v(751)
    assign n9186 = rst ? encrypted_data_buf[477] : encrypted_data_buf_next[477];   // modexp_top.v(751)
    assign n9187 = rst ? encrypted_data_buf[476] : encrypted_data_buf_next[476];   // modexp_top.v(751)
    assign n9188 = rst ? encrypted_data_buf[475] : encrypted_data_buf_next[475];   // modexp_top.v(751)
    assign n9189 = rst ? encrypted_data_buf[474] : encrypted_data_buf_next[474];   // modexp_top.v(751)
    assign n9190 = rst ? encrypted_data_buf[473] : encrypted_data_buf_next[473];   // modexp_top.v(751)
    assign n9191 = rst ? encrypted_data_buf[472] : encrypted_data_buf_next[472];   // modexp_top.v(751)
    assign n9192 = rst ? encrypted_data_buf[471] : encrypted_data_buf_next[471];   // modexp_top.v(751)
    assign n9193 = rst ? encrypted_data_buf[470] : encrypted_data_buf_next[470];   // modexp_top.v(751)
    assign n9194 = rst ? encrypted_data_buf[469] : encrypted_data_buf_next[469];   // modexp_top.v(751)
    assign n9195 = rst ? encrypted_data_buf[468] : encrypted_data_buf_next[468];   // modexp_top.v(751)
    assign n9196 = rst ? encrypted_data_buf[467] : encrypted_data_buf_next[467];   // modexp_top.v(751)
    assign n9197 = rst ? encrypted_data_buf[466] : encrypted_data_buf_next[466];   // modexp_top.v(751)
    assign n9198 = rst ? encrypted_data_buf[465] : encrypted_data_buf_next[465];   // modexp_top.v(751)
    assign n9199 = rst ? encrypted_data_buf[464] : encrypted_data_buf_next[464];   // modexp_top.v(751)
    assign n9200 = rst ? encrypted_data_buf[463] : encrypted_data_buf_next[463];   // modexp_top.v(751)
    assign n9201 = rst ? encrypted_data_buf[462] : encrypted_data_buf_next[462];   // modexp_top.v(751)
    assign n9202 = rst ? encrypted_data_buf[461] : encrypted_data_buf_next[461];   // modexp_top.v(751)
    assign n9203 = rst ? encrypted_data_buf[460] : encrypted_data_buf_next[460];   // modexp_top.v(751)
    assign n9204 = rst ? encrypted_data_buf[459] : encrypted_data_buf_next[459];   // modexp_top.v(751)
    assign n9205 = rst ? encrypted_data_buf[458] : encrypted_data_buf_next[458];   // modexp_top.v(751)
    assign n9206 = rst ? encrypted_data_buf[457] : encrypted_data_buf_next[457];   // modexp_top.v(751)
    assign n9207 = rst ? encrypted_data_buf[456] : encrypted_data_buf_next[456];   // modexp_top.v(751)
    assign n9208 = rst ? encrypted_data_buf[455] : encrypted_data_buf_next[455];   // modexp_top.v(751)
    assign n9209 = rst ? encrypted_data_buf[454] : encrypted_data_buf_next[454];   // modexp_top.v(751)
    assign n9210 = rst ? encrypted_data_buf[453] : encrypted_data_buf_next[453];   // modexp_top.v(751)
    assign n9211 = rst ? encrypted_data_buf[452] : encrypted_data_buf_next[452];   // modexp_top.v(751)
    assign n9212 = rst ? encrypted_data_buf[451] : encrypted_data_buf_next[451];   // modexp_top.v(751)
    assign n9213 = rst ? encrypted_data_buf[450] : encrypted_data_buf_next[450];   // modexp_top.v(751)
    assign n9214 = rst ? encrypted_data_buf[449] : encrypted_data_buf_next[449];   // modexp_top.v(751)
    assign n9215 = rst ? encrypted_data_buf[448] : encrypted_data_buf_next[448];   // modexp_top.v(751)
    assign n9216 = rst ? encrypted_data_buf[447] : encrypted_data_buf_next[447];   // modexp_top.v(751)
    assign n9217 = rst ? encrypted_data_buf[446] : encrypted_data_buf_next[446];   // modexp_top.v(751)
    assign n9218 = rst ? encrypted_data_buf[445] : encrypted_data_buf_next[445];   // modexp_top.v(751)
    assign n9219 = rst ? encrypted_data_buf[444] : encrypted_data_buf_next[444];   // modexp_top.v(751)
    assign n9220 = rst ? encrypted_data_buf[443] : encrypted_data_buf_next[443];   // modexp_top.v(751)
    assign n9221 = rst ? encrypted_data_buf[442] : encrypted_data_buf_next[442];   // modexp_top.v(751)
    assign n9222 = rst ? encrypted_data_buf[441] : encrypted_data_buf_next[441];   // modexp_top.v(751)
    assign n9223 = rst ? encrypted_data_buf[440] : encrypted_data_buf_next[440];   // modexp_top.v(751)
    assign n9224 = rst ? encrypted_data_buf[439] : encrypted_data_buf_next[439];   // modexp_top.v(751)
    assign n9225 = rst ? encrypted_data_buf[438] : encrypted_data_buf_next[438];   // modexp_top.v(751)
    assign n9226 = rst ? encrypted_data_buf[437] : encrypted_data_buf_next[437];   // modexp_top.v(751)
    assign n9227 = rst ? encrypted_data_buf[436] : encrypted_data_buf_next[436];   // modexp_top.v(751)
    assign n9228 = rst ? encrypted_data_buf[435] : encrypted_data_buf_next[435];   // modexp_top.v(751)
    assign n9229 = rst ? encrypted_data_buf[434] : encrypted_data_buf_next[434];   // modexp_top.v(751)
    assign n9230 = rst ? encrypted_data_buf[433] : encrypted_data_buf_next[433];   // modexp_top.v(751)
    assign n9231 = rst ? encrypted_data_buf[432] : encrypted_data_buf_next[432];   // modexp_top.v(751)
    assign n9232 = rst ? encrypted_data_buf[431] : encrypted_data_buf_next[431];   // modexp_top.v(751)
    assign n9233 = rst ? encrypted_data_buf[430] : encrypted_data_buf_next[430];   // modexp_top.v(751)
    assign n9234 = rst ? encrypted_data_buf[429] : encrypted_data_buf_next[429];   // modexp_top.v(751)
    assign n9235 = rst ? encrypted_data_buf[428] : encrypted_data_buf_next[428];   // modexp_top.v(751)
    assign n9236 = rst ? encrypted_data_buf[427] : encrypted_data_buf_next[427];   // modexp_top.v(751)
    assign n9237 = rst ? encrypted_data_buf[426] : encrypted_data_buf_next[426];   // modexp_top.v(751)
    assign n9238 = rst ? encrypted_data_buf[425] : encrypted_data_buf_next[425];   // modexp_top.v(751)
    assign n9239 = rst ? encrypted_data_buf[424] : encrypted_data_buf_next[424];   // modexp_top.v(751)
    assign n9240 = rst ? encrypted_data_buf[423] : encrypted_data_buf_next[423];   // modexp_top.v(751)
    assign n9241 = rst ? encrypted_data_buf[422] : encrypted_data_buf_next[422];   // modexp_top.v(751)
    assign n9242 = rst ? encrypted_data_buf[421] : encrypted_data_buf_next[421];   // modexp_top.v(751)
    assign n9243 = rst ? encrypted_data_buf[420] : encrypted_data_buf_next[420];   // modexp_top.v(751)
    assign n9244 = rst ? encrypted_data_buf[419] : encrypted_data_buf_next[419];   // modexp_top.v(751)
    assign n9245 = rst ? encrypted_data_buf[418] : encrypted_data_buf_next[418];   // modexp_top.v(751)
    assign n9246 = rst ? encrypted_data_buf[417] : encrypted_data_buf_next[417];   // modexp_top.v(751)
    assign n9247 = rst ? encrypted_data_buf[416] : encrypted_data_buf_next[416];   // modexp_top.v(751)
    assign n9248 = rst ? encrypted_data_buf[415] : encrypted_data_buf_next[415];   // modexp_top.v(751)
    assign n9249 = rst ? encrypted_data_buf[414] : encrypted_data_buf_next[414];   // modexp_top.v(751)
    assign n9250 = rst ? encrypted_data_buf[413] : encrypted_data_buf_next[413];   // modexp_top.v(751)
    assign n9251 = rst ? encrypted_data_buf[412] : encrypted_data_buf_next[412];   // modexp_top.v(751)
    assign n9252 = rst ? encrypted_data_buf[411] : encrypted_data_buf_next[411];   // modexp_top.v(751)
    assign n9253 = rst ? encrypted_data_buf[410] : encrypted_data_buf_next[410];   // modexp_top.v(751)
    assign n9254 = rst ? encrypted_data_buf[409] : encrypted_data_buf_next[409];   // modexp_top.v(751)
    assign n9255 = rst ? encrypted_data_buf[408] : encrypted_data_buf_next[408];   // modexp_top.v(751)
    assign n9256 = rst ? encrypted_data_buf[407] : encrypted_data_buf_next[407];   // modexp_top.v(751)
    assign n9257 = rst ? encrypted_data_buf[406] : encrypted_data_buf_next[406];   // modexp_top.v(751)
    assign n9258 = rst ? encrypted_data_buf[405] : encrypted_data_buf_next[405];   // modexp_top.v(751)
    assign n9259 = rst ? encrypted_data_buf[404] : encrypted_data_buf_next[404];   // modexp_top.v(751)
    assign n9260 = rst ? encrypted_data_buf[403] : encrypted_data_buf_next[403];   // modexp_top.v(751)
    assign n9261 = rst ? encrypted_data_buf[402] : encrypted_data_buf_next[402];   // modexp_top.v(751)
    assign n9262 = rst ? encrypted_data_buf[401] : encrypted_data_buf_next[401];   // modexp_top.v(751)
    assign n9263 = rst ? encrypted_data_buf[400] : encrypted_data_buf_next[400];   // modexp_top.v(751)
    assign n9264 = rst ? encrypted_data_buf[399] : encrypted_data_buf_next[399];   // modexp_top.v(751)
    assign n9265 = rst ? encrypted_data_buf[398] : encrypted_data_buf_next[398];   // modexp_top.v(751)
    assign n9266 = rst ? encrypted_data_buf[397] : encrypted_data_buf_next[397];   // modexp_top.v(751)
    assign n9267 = rst ? encrypted_data_buf[396] : encrypted_data_buf_next[396];   // modexp_top.v(751)
    assign n9268 = rst ? encrypted_data_buf[395] : encrypted_data_buf_next[395];   // modexp_top.v(751)
    assign n9269 = rst ? encrypted_data_buf[394] : encrypted_data_buf_next[394];   // modexp_top.v(751)
    assign n9270 = rst ? encrypted_data_buf[393] : encrypted_data_buf_next[393];   // modexp_top.v(751)
    assign n9271 = rst ? encrypted_data_buf[392] : encrypted_data_buf_next[392];   // modexp_top.v(751)
    assign n9272 = rst ? encrypted_data_buf[391] : encrypted_data_buf_next[391];   // modexp_top.v(751)
    assign n9273 = rst ? encrypted_data_buf[390] : encrypted_data_buf_next[390];   // modexp_top.v(751)
    assign n9274 = rst ? encrypted_data_buf[389] : encrypted_data_buf_next[389];   // modexp_top.v(751)
    assign n9275 = rst ? encrypted_data_buf[388] : encrypted_data_buf_next[388];   // modexp_top.v(751)
    assign n9276 = rst ? encrypted_data_buf[387] : encrypted_data_buf_next[387];   // modexp_top.v(751)
    assign n9277 = rst ? encrypted_data_buf[386] : encrypted_data_buf_next[386];   // modexp_top.v(751)
    assign n9278 = rst ? encrypted_data_buf[385] : encrypted_data_buf_next[385];   // modexp_top.v(751)
    assign n9279 = rst ? encrypted_data_buf[384] : encrypted_data_buf_next[384];   // modexp_top.v(751)
    assign n9280 = rst ? encrypted_data_buf[383] : encrypted_data_buf_next[383];   // modexp_top.v(751)
    assign n9281 = rst ? encrypted_data_buf[382] : encrypted_data_buf_next[382];   // modexp_top.v(751)
    assign n9282 = rst ? encrypted_data_buf[381] : encrypted_data_buf_next[381];   // modexp_top.v(751)
    assign n9283 = rst ? encrypted_data_buf[380] : encrypted_data_buf_next[380];   // modexp_top.v(751)
    assign n9284 = rst ? encrypted_data_buf[379] : encrypted_data_buf_next[379];   // modexp_top.v(751)
    assign n9285 = rst ? encrypted_data_buf[378] : encrypted_data_buf_next[378];   // modexp_top.v(751)
    assign n9286 = rst ? encrypted_data_buf[377] : encrypted_data_buf_next[377];   // modexp_top.v(751)
    assign n9287 = rst ? encrypted_data_buf[376] : encrypted_data_buf_next[376];   // modexp_top.v(751)
    assign n9288 = rst ? encrypted_data_buf[375] : encrypted_data_buf_next[375];   // modexp_top.v(751)
    assign n9289 = rst ? encrypted_data_buf[374] : encrypted_data_buf_next[374];   // modexp_top.v(751)
    assign n9290 = rst ? encrypted_data_buf[373] : encrypted_data_buf_next[373];   // modexp_top.v(751)
    assign n9291 = rst ? encrypted_data_buf[372] : encrypted_data_buf_next[372];   // modexp_top.v(751)
    assign n9292 = rst ? encrypted_data_buf[371] : encrypted_data_buf_next[371];   // modexp_top.v(751)
    assign n9293 = rst ? encrypted_data_buf[370] : encrypted_data_buf_next[370];   // modexp_top.v(751)
    assign n9294 = rst ? encrypted_data_buf[369] : encrypted_data_buf_next[369];   // modexp_top.v(751)
    assign n9295 = rst ? encrypted_data_buf[368] : encrypted_data_buf_next[368];   // modexp_top.v(751)
    assign n9296 = rst ? encrypted_data_buf[367] : encrypted_data_buf_next[367];   // modexp_top.v(751)
    assign n9297 = rst ? encrypted_data_buf[366] : encrypted_data_buf_next[366];   // modexp_top.v(751)
    assign n9298 = rst ? encrypted_data_buf[365] : encrypted_data_buf_next[365];   // modexp_top.v(751)
    assign n9299 = rst ? encrypted_data_buf[364] : encrypted_data_buf_next[364];   // modexp_top.v(751)
    assign n9300 = rst ? encrypted_data_buf[363] : encrypted_data_buf_next[363];   // modexp_top.v(751)
    assign n9301 = rst ? encrypted_data_buf[362] : encrypted_data_buf_next[362];   // modexp_top.v(751)
    assign n9302 = rst ? encrypted_data_buf[361] : encrypted_data_buf_next[361];   // modexp_top.v(751)
    assign n9303 = rst ? encrypted_data_buf[360] : encrypted_data_buf_next[360];   // modexp_top.v(751)
    assign n9304 = rst ? encrypted_data_buf[359] : encrypted_data_buf_next[359];   // modexp_top.v(751)
    assign n9305 = rst ? encrypted_data_buf[358] : encrypted_data_buf_next[358];   // modexp_top.v(751)
    assign n9306 = rst ? encrypted_data_buf[357] : encrypted_data_buf_next[357];   // modexp_top.v(751)
    assign n9307 = rst ? encrypted_data_buf[356] : encrypted_data_buf_next[356];   // modexp_top.v(751)
    assign n9308 = rst ? encrypted_data_buf[355] : encrypted_data_buf_next[355];   // modexp_top.v(751)
    assign n9309 = rst ? encrypted_data_buf[354] : encrypted_data_buf_next[354];   // modexp_top.v(751)
    assign n9310 = rst ? encrypted_data_buf[353] : encrypted_data_buf_next[353];   // modexp_top.v(751)
    assign n9311 = rst ? encrypted_data_buf[352] : encrypted_data_buf_next[352];   // modexp_top.v(751)
    assign n9312 = rst ? encrypted_data_buf[351] : encrypted_data_buf_next[351];   // modexp_top.v(751)
    assign n9313 = rst ? encrypted_data_buf[350] : encrypted_data_buf_next[350];   // modexp_top.v(751)
    assign n9314 = rst ? encrypted_data_buf[349] : encrypted_data_buf_next[349];   // modexp_top.v(751)
    assign n9315 = rst ? encrypted_data_buf[348] : encrypted_data_buf_next[348];   // modexp_top.v(751)
    assign n9316 = rst ? encrypted_data_buf[347] : encrypted_data_buf_next[347];   // modexp_top.v(751)
    assign n9317 = rst ? encrypted_data_buf[346] : encrypted_data_buf_next[346];   // modexp_top.v(751)
    assign n9318 = rst ? encrypted_data_buf[345] : encrypted_data_buf_next[345];   // modexp_top.v(751)
    assign n9319 = rst ? encrypted_data_buf[344] : encrypted_data_buf_next[344];   // modexp_top.v(751)
    assign n9320 = rst ? encrypted_data_buf[343] : encrypted_data_buf_next[343];   // modexp_top.v(751)
    assign n9321 = rst ? encrypted_data_buf[342] : encrypted_data_buf_next[342];   // modexp_top.v(751)
    assign n9322 = rst ? encrypted_data_buf[341] : encrypted_data_buf_next[341];   // modexp_top.v(751)
    assign n9323 = rst ? encrypted_data_buf[340] : encrypted_data_buf_next[340];   // modexp_top.v(751)
    assign n9324 = rst ? encrypted_data_buf[339] : encrypted_data_buf_next[339];   // modexp_top.v(751)
    assign n9325 = rst ? encrypted_data_buf[338] : encrypted_data_buf_next[338];   // modexp_top.v(751)
    assign n9326 = rst ? encrypted_data_buf[337] : encrypted_data_buf_next[337];   // modexp_top.v(751)
    assign n9327 = rst ? encrypted_data_buf[336] : encrypted_data_buf_next[336];   // modexp_top.v(751)
    assign n9328 = rst ? encrypted_data_buf[335] : encrypted_data_buf_next[335];   // modexp_top.v(751)
    assign n9329 = rst ? encrypted_data_buf[334] : encrypted_data_buf_next[334];   // modexp_top.v(751)
    assign n9330 = rst ? encrypted_data_buf[333] : encrypted_data_buf_next[333];   // modexp_top.v(751)
    assign n9331 = rst ? encrypted_data_buf[332] : encrypted_data_buf_next[332];   // modexp_top.v(751)
    assign n9332 = rst ? encrypted_data_buf[331] : encrypted_data_buf_next[331];   // modexp_top.v(751)
    assign n9333 = rst ? encrypted_data_buf[330] : encrypted_data_buf_next[330];   // modexp_top.v(751)
    assign n9334 = rst ? encrypted_data_buf[329] : encrypted_data_buf_next[329];   // modexp_top.v(751)
    assign n9335 = rst ? encrypted_data_buf[328] : encrypted_data_buf_next[328];   // modexp_top.v(751)
    assign n9336 = rst ? encrypted_data_buf[327] : encrypted_data_buf_next[327];   // modexp_top.v(751)
    assign n9337 = rst ? encrypted_data_buf[326] : encrypted_data_buf_next[326];   // modexp_top.v(751)
    assign n9338 = rst ? encrypted_data_buf[325] : encrypted_data_buf_next[325];   // modexp_top.v(751)
    assign n9339 = rst ? encrypted_data_buf[324] : encrypted_data_buf_next[324];   // modexp_top.v(751)
    assign n9340 = rst ? encrypted_data_buf[323] : encrypted_data_buf_next[323];   // modexp_top.v(751)
    assign n9341 = rst ? encrypted_data_buf[322] : encrypted_data_buf_next[322];   // modexp_top.v(751)
    assign n9342 = rst ? encrypted_data_buf[321] : encrypted_data_buf_next[321];   // modexp_top.v(751)
    assign n9343 = rst ? encrypted_data_buf[320] : encrypted_data_buf_next[320];   // modexp_top.v(751)
    assign n9344 = rst ? encrypted_data_buf[319] : encrypted_data_buf_next[319];   // modexp_top.v(751)
    assign n9345 = rst ? encrypted_data_buf[318] : encrypted_data_buf_next[318];   // modexp_top.v(751)
    assign n9346 = rst ? encrypted_data_buf[317] : encrypted_data_buf_next[317];   // modexp_top.v(751)
    assign n9347 = rst ? encrypted_data_buf[316] : encrypted_data_buf_next[316];   // modexp_top.v(751)
    assign n9348 = rst ? encrypted_data_buf[315] : encrypted_data_buf_next[315];   // modexp_top.v(751)
    assign n9349 = rst ? encrypted_data_buf[314] : encrypted_data_buf_next[314];   // modexp_top.v(751)
    assign n9350 = rst ? encrypted_data_buf[313] : encrypted_data_buf_next[313];   // modexp_top.v(751)
    assign n9351 = rst ? encrypted_data_buf[312] : encrypted_data_buf_next[312];   // modexp_top.v(751)
    assign n9352 = rst ? encrypted_data_buf[311] : encrypted_data_buf_next[311];   // modexp_top.v(751)
    assign n9353 = rst ? encrypted_data_buf[310] : encrypted_data_buf_next[310];   // modexp_top.v(751)
    assign n9354 = rst ? encrypted_data_buf[309] : encrypted_data_buf_next[309];   // modexp_top.v(751)
    assign n9355 = rst ? encrypted_data_buf[308] : encrypted_data_buf_next[308];   // modexp_top.v(751)
    assign n9356 = rst ? encrypted_data_buf[307] : encrypted_data_buf_next[307];   // modexp_top.v(751)
    assign n9357 = rst ? encrypted_data_buf[306] : encrypted_data_buf_next[306];   // modexp_top.v(751)
    assign n9358 = rst ? encrypted_data_buf[305] : encrypted_data_buf_next[305];   // modexp_top.v(751)
    assign n9359 = rst ? encrypted_data_buf[304] : encrypted_data_buf_next[304];   // modexp_top.v(751)
    assign n9360 = rst ? encrypted_data_buf[303] : encrypted_data_buf_next[303];   // modexp_top.v(751)
    assign n9361 = rst ? encrypted_data_buf[302] : encrypted_data_buf_next[302];   // modexp_top.v(751)
    assign n9362 = rst ? encrypted_data_buf[301] : encrypted_data_buf_next[301];   // modexp_top.v(751)
    assign n9363 = rst ? encrypted_data_buf[300] : encrypted_data_buf_next[300];   // modexp_top.v(751)
    assign n9364 = rst ? encrypted_data_buf[299] : encrypted_data_buf_next[299];   // modexp_top.v(751)
    assign n9365 = rst ? encrypted_data_buf[298] : encrypted_data_buf_next[298];   // modexp_top.v(751)
    assign n9366 = rst ? encrypted_data_buf[297] : encrypted_data_buf_next[297];   // modexp_top.v(751)
    assign n9367 = rst ? encrypted_data_buf[296] : encrypted_data_buf_next[296];   // modexp_top.v(751)
    assign n9368 = rst ? encrypted_data_buf[295] : encrypted_data_buf_next[295];   // modexp_top.v(751)
    assign n9369 = rst ? encrypted_data_buf[294] : encrypted_data_buf_next[294];   // modexp_top.v(751)
    assign n9370 = rst ? encrypted_data_buf[293] : encrypted_data_buf_next[293];   // modexp_top.v(751)
    assign n9371 = rst ? encrypted_data_buf[292] : encrypted_data_buf_next[292];   // modexp_top.v(751)
    assign n9372 = rst ? encrypted_data_buf[291] : encrypted_data_buf_next[291];   // modexp_top.v(751)
    assign n9373 = rst ? encrypted_data_buf[290] : encrypted_data_buf_next[290];   // modexp_top.v(751)
    assign n9374 = rst ? encrypted_data_buf[289] : encrypted_data_buf_next[289];   // modexp_top.v(751)
    assign n9375 = rst ? encrypted_data_buf[288] : encrypted_data_buf_next[288];   // modexp_top.v(751)
    assign n9376 = rst ? encrypted_data_buf[287] : encrypted_data_buf_next[287];   // modexp_top.v(751)
    assign n9377 = rst ? encrypted_data_buf[286] : encrypted_data_buf_next[286];   // modexp_top.v(751)
    assign n9378 = rst ? encrypted_data_buf[285] : encrypted_data_buf_next[285];   // modexp_top.v(751)
    assign n9379 = rst ? encrypted_data_buf[284] : encrypted_data_buf_next[284];   // modexp_top.v(751)
    assign n9380 = rst ? encrypted_data_buf[283] : encrypted_data_buf_next[283];   // modexp_top.v(751)
    assign n9381 = rst ? encrypted_data_buf[282] : encrypted_data_buf_next[282];   // modexp_top.v(751)
    assign n9382 = rst ? encrypted_data_buf[281] : encrypted_data_buf_next[281];   // modexp_top.v(751)
    assign n9383 = rst ? encrypted_data_buf[280] : encrypted_data_buf_next[280];   // modexp_top.v(751)
    assign n9384 = rst ? encrypted_data_buf[279] : encrypted_data_buf_next[279];   // modexp_top.v(751)
    assign n9385 = rst ? encrypted_data_buf[278] : encrypted_data_buf_next[278];   // modexp_top.v(751)
    assign n9386 = rst ? encrypted_data_buf[277] : encrypted_data_buf_next[277];   // modexp_top.v(751)
    assign n9387 = rst ? encrypted_data_buf[276] : encrypted_data_buf_next[276];   // modexp_top.v(751)
    assign n9388 = rst ? encrypted_data_buf[275] : encrypted_data_buf_next[275];   // modexp_top.v(751)
    assign n9389 = rst ? encrypted_data_buf[274] : encrypted_data_buf_next[274];   // modexp_top.v(751)
    assign n9390 = rst ? encrypted_data_buf[273] : encrypted_data_buf_next[273];   // modexp_top.v(751)
    assign n9391 = rst ? encrypted_data_buf[272] : encrypted_data_buf_next[272];   // modexp_top.v(751)
    assign n9392 = rst ? encrypted_data_buf[271] : encrypted_data_buf_next[271];   // modexp_top.v(751)
    assign n9393 = rst ? encrypted_data_buf[270] : encrypted_data_buf_next[270];   // modexp_top.v(751)
    assign n9394 = rst ? encrypted_data_buf[269] : encrypted_data_buf_next[269];   // modexp_top.v(751)
    assign n9395 = rst ? encrypted_data_buf[268] : encrypted_data_buf_next[268];   // modexp_top.v(751)
    assign n9396 = rst ? encrypted_data_buf[267] : encrypted_data_buf_next[267];   // modexp_top.v(751)
    assign n9397 = rst ? encrypted_data_buf[266] : encrypted_data_buf_next[266];   // modexp_top.v(751)
    assign n9398 = rst ? encrypted_data_buf[265] : encrypted_data_buf_next[265];   // modexp_top.v(751)
    assign n9399 = rst ? encrypted_data_buf[264] : encrypted_data_buf_next[264];   // modexp_top.v(751)
    assign n9400 = rst ? encrypted_data_buf[263] : encrypted_data_buf_next[263];   // modexp_top.v(751)
    assign n9401 = rst ? encrypted_data_buf[262] : encrypted_data_buf_next[262];   // modexp_top.v(751)
    assign n9402 = rst ? encrypted_data_buf[261] : encrypted_data_buf_next[261];   // modexp_top.v(751)
    assign n9403 = rst ? encrypted_data_buf[260] : encrypted_data_buf_next[260];   // modexp_top.v(751)
    assign n9404 = rst ? encrypted_data_buf[259] : encrypted_data_buf_next[259];   // modexp_top.v(751)
    assign n9405 = rst ? encrypted_data_buf[258] : encrypted_data_buf_next[258];   // modexp_top.v(751)
    assign n9406 = rst ? encrypted_data_buf[257] : encrypted_data_buf_next[257];   // modexp_top.v(751)
    assign n9407 = rst ? encrypted_data_buf[256] : encrypted_data_buf_next[256];   // modexp_top.v(751)
    assign n9408 = rst ? encrypted_data_buf[255] : encrypted_data_buf_next[255];   // modexp_top.v(751)
    assign n9409 = rst ? encrypted_data_buf[254] : encrypted_data_buf_next[254];   // modexp_top.v(751)
    assign n9410 = rst ? encrypted_data_buf[253] : encrypted_data_buf_next[253];   // modexp_top.v(751)
    assign n9411 = rst ? encrypted_data_buf[252] : encrypted_data_buf_next[252];   // modexp_top.v(751)
    assign n9412 = rst ? encrypted_data_buf[251] : encrypted_data_buf_next[251];   // modexp_top.v(751)
    assign n9413 = rst ? encrypted_data_buf[250] : encrypted_data_buf_next[250];   // modexp_top.v(751)
    assign n9414 = rst ? encrypted_data_buf[249] : encrypted_data_buf_next[249];   // modexp_top.v(751)
    assign n9415 = rst ? encrypted_data_buf[248] : encrypted_data_buf_next[248];   // modexp_top.v(751)
    assign n9416 = rst ? encrypted_data_buf[247] : encrypted_data_buf_next[247];   // modexp_top.v(751)
    assign n9417 = rst ? encrypted_data_buf[246] : encrypted_data_buf_next[246];   // modexp_top.v(751)
    assign n9418 = rst ? encrypted_data_buf[245] : encrypted_data_buf_next[245];   // modexp_top.v(751)
    assign n9419 = rst ? encrypted_data_buf[244] : encrypted_data_buf_next[244];   // modexp_top.v(751)
    assign n9420 = rst ? encrypted_data_buf[243] : encrypted_data_buf_next[243];   // modexp_top.v(751)
    assign n9421 = rst ? encrypted_data_buf[242] : encrypted_data_buf_next[242];   // modexp_top.v(751)
    assign n9422 = rst ? encrypted_data_buf[241] : encrypted_data_buf_next[241];   // modexp_top.v(751)
    assign n9423 = rst ? encrypted_data_buf[240] : encrypted_data_buf_next[240];   // modexp_top.v(751)
    assign n9424 = rst ? encrypted_data_buf[239] : encrypted_data_buf_next[239];   // modexp_top.v(751)
    assign n9425 = rst ? encrypted_data_buf[238] : encrypted_data_buf_next[238];   // modexp_top.v(751)
    assign n9426 = rst ? encrypted_data_buf[237] : encrypted_data_buf_next[237];   // modexp_top.v(751)
    assign n9427 = rst ? encrypted_data_buf[236] : encrypted_data_buf_next[236];   // modexp_top.v(751)
    assign n9428 = rst ? encrypted_data_buf[235] : encrypted_data_buf_next[235];   // modexp_top.v(751)
    assign n9429 = rst ? encrypted_data_buf[234] : encrypted_data_buf_next[234];   // modexp_top.v(751)
    assign n9430 = rst ? encrypted_data_buf[233] : encrypted_data_buf_next[233];   // modexp_top.v(751)
    assign n9431 = rst ? encrypted_data_buf[232] : encrypted_data_buf_next[232];   // modexp_top.v(751)
    assign n9432 = rst ? encrypted_data_buf[231] : encrypted_data_buf_next[231];   // modexp_top.v(751)
    assign n9433 = rst ? encrypted_data_buf[230] : encrypted_data_buf_next[230];   // modexp_top.v(751)
    assign n9434 = rst ? encrypted_data_buf[229] : encrypted_data_buf_next[229];   // modexp_top.v(751)
    assign n9435 = rst ? encrypted_data_buf[228] : encrypted_data_buf_next[228];   // modexp_top.v(751)
    assign n9436 = rst ? encrypted_data_buf[227] : encrypted_data_buf_next[227];   // modexp_top.v(751)
    assign n9437 = rst ? encrypted_data_buf[226] : encrypted_data_buf_next[226];   // modexp_top.v(751)
    assign n9438 = rst ? encrypted_data_buf[225] : encrypted_data_buf_next[225];   // modexp_top.v(751)
    assign n9439 = rst ? encrypted_data_buf[224] : encrypted_data_buf_next[224];   // modexp_top.v(751)
    assign n9440 = rst ? encrypted_data_buf[223] : encrypted_data_buf_next[223];   // modexp_top.v(751)
    assign n9441 = rst ? encrypted_data_buf[222] : encrypted_data_buf_next[222];   // modexp_top.v(751)
    assign n9442 = rst ? encrypted_data_buf[221] : encrypted_data_buf_next[221];   // modexp_top.v(751)
    assign n9443 = rst ? encrypted_data_buf[220] : encrypted_data_buf_next[220];   // modexp_top.v(751)
    assign n9444 = rst ? encrypted_data_buf[219] : encrypted_data_buf_next[219];   // modexp_top.v(751)
    assign n9445 = rst ? encrypted_data_buf[218] : encrypted_data_buf_next[218];   // modexp_top.v(751)
    assign n9446 = rst ? encrypted_data_buf[217] : encrypted_data_buf_next[217];   // modexp_top.v(751)
    assign n9447 = rst ? encrypted_data_buf[216] : encrypted_data_buf_next[216];   // modexp_top.v(751)
    assign n9448 = rst ? encrypted_data_buf[215] : encrypted_data_buf_next[215];   // modexp_top.v(751)
    assign n9449 = rst ? encrypted_data_buf[214] : encrypted_data_buf_next[214];   // modexp_top.v(751)
    assign n9450 = rst ? encrypted_data_buf[213] : encrypted_data_buf_next[213];   // modexp_top.v(751)
    assign n9451 = rst ? encrypted_data_buf[212] : encrypted_data_buf_next[212];   // modexp_top.v(751)
    assign n9452 = rst ? encrypted_data_buf[211] : encrypted_data_buf_next[211];   // modexp_top.v(751)
    assign n9453 = rst ? encrypted_data_buf[210] : encrypted_data_buf_next[210];   // modexp_top.v(751)
    assign n9454 = rst ? encrypted_data_buf[209] : encrypted_data_buf_next[209];   // modexp_top.v(751)
    assign n9455 = rst ? encrypted_data_buf[208] : encrypted_data_buf_next[208];   // modexp_top.v(751)
    assign n9456 = rst ? encrypted_data_buf[207] : encrypted_data_buf_next[207];   // modexp_top.v(751)
    assign n9457 = rst ? encrypted_data_buf[206] : encrypted_data_buf_next[206];   // modexp_top.v(751)
    assign n9458 = rst ? encrypted_data_buf[205] : encrypted_data_buf_next[205];   // modexp_top.v(751)
    assign n9459 = rst ? encrypted_data_buf[204] : encrypted_data_buf_next[204];   // modexp_top.v(751)
    assign n9460 = rst ? encrypted_data_buf[203] : encrypted_data_buf_next[203];   // modexp_top.v(751)
    assign n9461 = rst ? encrypted_data_buf[202] : encrypted_data_buf_next[202];   // modexp_top.v(751)
    assign n9462 = rst ? encrypted_data_buf[201] : encrypted_data_buf_next[201];   // modexp_top.v(751)
    assign n9463 = rst ? encrypted_data_buf[200] : encrypted_data_buf_next[200];   // modexp_top.v(751)
    assign n9464 = rst ? encrypted_data_buf[199] : encrypted_data_buf_next[199];   // modexp_top.v(751)
    assign n9465 = rst ? encrypted_data_buf[198] : encrypted_data_buf_next[198];   // modexp_top.v(751)
    assign n9466 = rst ? encrypted_data_buf[197] : encrypted_data_buf_next[197];   // modexp_top.v(751)
    assign n9467 = rst ? encrypted_data_buf[196] : encrypted_data_buf_next[196];   // modexp_top.v(751)
    assign n9468 = rst ? encrypted_data_buf[195] : encrypted_data_buf_next[195];   // modexp_top.v(751)
    assign n9469 = rst ? encrypted_data_buf[194] : encrypted_data_buf_next[194];   // modexp_top.v(751)
    assign n9470 = rst ? encrypted_data_buf[193] : encrypted_data_buf_next[193];   // modexp_top.v(751)
    assign n9471 = rst ? encrypted_data_buf[192] : encrypted_data_buf_next[192];   // modexp_top.v(751)
    assign n9472 = rst ? encrypted_data_buf[191] : encrypted_data_buf_next[191];   // modexp_top.v(751)
    assign n9473 = rst ? encrypted_data_buf[190] : encrypted_data_buf_next[190];   // modexp_top.v(751)
    assign n9474 = rst ? encrypted_data_buf[189] : encrypted_data_buf_next[189];   // modexp_top.v(751)
    assign n9475 = rst ? encrypted_data_buf[188] : encrypted_data_buf_next[188];   // modexp_top.v(751)
    assign n9476 = rst ? encrypted_data_buf[187] : encrypted_data_buf_next[187];   // modexp_top.v(751)
    assign n9477 = rst ? encrypted_data_buf[186] : encrypted_data_buf_next[186];   // modexp_top.v(751)
    assign n9478 = rst ? encrypted_data_buf[185] : encrypted_data_buf_next[185];   // modexp_top.v(751)
    assign n9479 = rst ? encrypted_data_buf[184] : encrypted_data_buf_next[184];   // modexp_top.v(751)
    assign n9480 = rst ? encrypted_data_buf[183] : encrypted_data_buf_next[183];   // modexp_top.v(751)
    assign n9481 = rst ? encrypted_data_buf[182] : encrypted_data_buf_next[182];   // modexp_top.v(751)
    assign n9482 = rst ? encrypted_data_buf[181] : encrypted_data_buf_next[181];   // modexp_top.v(751)
    assign n9483 = rst ? encrypted_data_buf[180] : encrypted_data_buf_next[180];   // modexp_top.v(751)
    assign n9484 = rst ? encrypted_data_buf[179] : encrypted_data_buf_next[179];   // modexp_top.v(751)
    assign n9485 = rst ? encrypted_data_buf[178] : encrypted_data_buf_next[178];   // modexp_top.v(751)
    assign n9486 = rst ? encrypted_data_buf[177] : encrypted_data_buf_next[177];   // modexp_top.v(751)
    assign n9487 = rst ? encrypted_data_buf[176] : encrypted_data_buf_next[176];   // modexp_top.v(751)
    assign n9488 = rst ? encrypted_data_buf[175] : encrypted_data_buf_next[175];   // modexp_top.v(751)
    assign n9489 = rst ? encrypted_data_buf[174] : encrypted_data_buf_next[174];   // modexp_top.v(751)
    assign n9490 = rst ? encrypted_data_buf[173] : encrypted_data_buf_next[173];   // modexp_top.v(751)
    assign n9491 = rst ? encrypted_data_buf[172] : encrypted_data_buf_next[172];   // modexp_top.v(751)
    assign n9492 = rst ? encrypted_data_buf[171] : encrypted_data_buf_next[171];   // modexp_top.v(751)
    assign n9493 = rst ? encrypted_data_buf[170] : encrypted_data_buf_next[170];   // modexp_top.v(751)
    assign n9494 = rst ? encrypted_data_buf[169] : encrypted_data_buf_next[169];   // modexp_top.v(751)
    assign n9495 = rst ? encrypted_data_buf[168] : encrypted_data_buf_next[168];   // modexp_top.v(751)
    assign n9496 = rst ? encrypted_data_buf[167] : encrypted_data_buf_next[167];   // modexp_top.v(751)
    assign n9497 = rst ? encrypted_data_buf[166] : encrypted_data_buf_next[166];   // modexp_top.v(751)
    assign n9498 = rst ? encrypted_data_buf[165] : encrypted_data_buf_next[165];   // modexp_top.v(751)
    assign n9499 = rst ? encrypted_data_buf[164] : encrypted_data_buf_next[164];   // modexp_top.v(751)
    assign n9500 = rst ? encrypted_data_buf[163] : encrypted_data_buf_next[163];   // modexp_top.v(751)
    assign n9501 = rst ? encrypted_data_buf[162] : encrypted_data_buf_next[162];   // modexp_top.v(751)
    assign n9502 = rst ? encrypted_data_buf[161] : encrypted_data_buf_next[161];   // modexp_top.v(751)
    assign n9503 = rst ? encrypted_data_buf[160] : encrypted_data_buf_next[160];   // modexp_top.v(751)
    assign n9504 = rst ? encrypted_data_buf[159] : encrypted_data_buf_next[159];   // modexp_top.v(751)
    assign n9505 = rst ? encrypted_data_buf[158] : encrypted_data_buf_next[158];   // modexp_top.v(751)
    assign n9506 = rst ? encrypted_data_buf[157] : encrypted_data_buf_next[157];   // modexp_top.v(751)
    assign n9507 = rst ? encrypted_data_buf[156] : encrypted_data_buf_next[156];   // modexp_top.v(751)
    assign n9508 = rst ? encrypted_data_buf[155] : encrypted_data_buf_next[155];   // modexp_top.v(751)
    assign n9509 = rst ? encrypted_data_buf[154] : encrypted_data_buf_next[154];   // modexp_top.v(751)
    assign n9510 = rst ? encrypted_data_buf[153] : encrypted_data_buf_next[153];   // modexp_top.v(751)
    assign n9511 = rst ? encrypted_data_buf[152] : encrypted_data_buf_next[152];   // modexp_top.v(751)
    assign n9512 = rst ? encrypted_data_buf[151] : encrypted_data_buf_next[151];   // modexp_top.v(751)
    assign n9513 = rst ? encrypted_data_buf[150] : encrypted_data_buf_next[150];   // modexp_top.v(751)
    assign n9514 = rst ? encrypted_data_buf[149] : encrypted_data_buf_next[149];   // modexp_top.v(751)
    assign n9515 = rst ? encrypted_data_buf[148] : encrypted_data_buf_next[148];   // modexp_top.v(751)
    assign n9516 = rst ? encrypted_data_buf[147] : encrypted_data_buf_next[147];   // modexp_top.v(751)
    assign n9517 = rst ? encrypted_data_buf[146] : encrypted_data_buf_next[146];   // modexp_top.v(751)
    assign n9518 = rst ? encrypted_data_buf[145] : encrypted_data_buf_next[145];   // modexp_top.v(751)
    assign n9519 = rst ? encrypted_data_buf[144] : encrypted_data_buf_next[144];   // modexp_top.v(751)
    assign n9520 = rst ? encrypted_data_buf[143] : encrypted_data_buf_next[143];   // modexp_top.v(751)
    assign n9521 = rst ? encrypted_data_buf[142] : encrypted_data_buf_next[142];   // modexp_top.v(751)
    assign n9522 = rst ? encrypted_data_buf[141] : encrypted_data_buf_next[141];   // modexp_top.v(751)
    assign n9523 = rst ? encrypted_data_buf[140] : encrypted_data_buf_next[140];   // modexp_top.v(751)
    assign n9524 = rst ? encrypted_data_buf[139] : encrypted_data_buf_next[139];   // modexp_top.v(751)
    assign n9525 = rst ? encrypted_data_buf[138] : encrypted_data_buf_next[138];   // modexp_top.v(751)
    assign n9526 = rst ? encrypted_data_buf[137] : encrypted_data_buf_next[137];   // modexp_top.v(751)
    assign n9527 = rst ? encrypted_data_buf[136] : encrypted_data_buf_next[136];   // modexp_top.v(751)
    assign n9528 = rst ? encrypted_data_buf[135] : encrypted_data_buf_next[135];   // modexp_top.v(751)
    assign n9529 = rst ? encrypted_data_buf[134] : encrypted_data_buf_next[134];   // modexp_top.v(751)
    assign n9530 = rst ? encrypted_data_buf[133] : encrypted_data_buf_next[133];   // modexp_top.v(751)
    assign n9531 = rst ? encrypted_data_buf[132] : encrypted_data_buf_next[132];   // modexp_top.v(751)
    assign n9532 = rst ? encrypted_data_buf[131] : encrypted_data_buf_next[131];   // modexp_top.v(751)
    assign n9533 = rst ? encrypted_data_buf[130] : encrypted_data_buf_next[130];   // modexp_top.v(751)
    assign n9534 = rst ? encrypted_data_buf[129] : encrypted_data_buf_next[129];   // modexp_top.v(751)
    assign n9535 = rst ? encrypted_data_buf[128] : encrypted_data_buf_next[128];   // modexp_top.v(751)
    assign n9536 = rst ? encrypted_data_buf[127] : encrypted_data_buf_next[127];   // modexp_top.v(751)
    assign n9537 = rst ? encrypted_data_buf[126] : encrypted_data_buf_next[126];   // modexp_top.v(751)
    assign n9538 = rst ? encrypted_data_buf[125] : encrypted_data_buf_next[125];   // modexp_top.v(751)
    assign n9539 = rst ? encrypted_data_buf[124] : encrypted_data_buf_next[124];   // modexp_top.v(751)
    assign n9540 = rst ? encrypted_data_buf[123] : encrypted_data_buf_next[123];   // modexp_top.v(751)
    assign n9541 = rst ? encrypted_data_buf[122] : encrypted_data_buf_next[122];   // modexp_top.v(751)
    assign n9542 = rst ? encrypted_data_buf[121] : encrypted_data_buf_next[121];   // modexp_top.v(751)
    assign n9543 = rst ? encrypted_data_buf[120] : encrypted_data_buf_next[120];   // modexp_top.v(751)
    assign n9544 = rst ? encrypted_data_buf[119] : encrypted_data_buf_next[119];   // modexp_top.v(751)
    assign n9545 = rst ? encrypted_data_buf[118] : encrypted_data_buf_next[118];   // modexp_top.v(751)
    assign n9546 = rst ? encrypted_data_buf[117] : encrypted_data_buf_next[117];   // modexp_top.v(751)
    assign n9547 = rst ? encrypted_data_buf[116] : encrypted_data_buf_next[116];   // modexp_top.v(751)
    assign n9548 = rst ? encrypted_data_buf[115] : encrypted_data_buf_next[115];   // modexp_top.v(751)
    assign n9549 = rst ? encrypted_data_buf[114] : encrypted_data_buf_next[114];   // modexp_top.v(751)
    assign n9550 = rst ? encrypted_data_buf[113] : encrypted_data_buf_next[113];   // modexp_top.v(751)
    assign n9551 = rst ? encrypted_data_buf[112] : encrypted_data_buf_next[112];   // modexp_top.v(751)
    assign n9552 = rst ? encrypted_data_buf[111] : encrypted_data_buf_next[111];   // modexp_top.v(751)
    assign n9553 = rst ? encrypted_data_buf[110] : encrypted_data_buf_next[110];   // modexp_top.v(751)
    assign n9554 = rst ? encrypted_data_buf[109] : encrypted_data_buf_next[109];   // modexp_top.v(751)
    assign n9555 = rst ? encrypted_data_buf[108] : encrypted_data_buf_next[108];   // modexp_top.v(751)
    assign n9556 = rst ? encrypted_data_buf[107] : encrypted_data_buf_next[107];   // modexp_top.v(751)
    assign n9557 = rst ? encrypted_data_buf[106] : encrypted_data_buf_next[106];   // modexp_top.v(751)
    assign n9558 = rst ? encrypted_data_buf[105] : encrypted_data_buf_next[105];   // modexp_top.v(751)
    assign n9559 = rst ? encrypted_data_buf[104] : encrypted_data_buf_next[104];   // modexp_top.v(751)
    assign n9560 = rst ? encrypted_data_buf[103] : encrypted_data_buf_next[103];   // modexp_top.v(751)
    assign n9561 = rst ? encrypted_data_buf[102] : encrypted_data_buf_next[102];   // modexp_top.v(751)
    assign n9562 = rst ? encrypted_data_buf[101] : encrypted_data_buf_next[101];   // modexp_top.v(751)
    assign n9563 = rst ? encrypted_data_buf[100] : encrypted_data_buf_next[100];   // modexp_top.v(751)
    assign n9564 = rst ? encrypted_data_buf[99] : encrypted_data_buf_next[99];   // modexp_top.v(751)
    assign n9565 = rst ? encrypted_data_buf[98] : encrypted_data_buf_next[98];   // modexp_top.v(751)
    assign n9566 = rst ? encrypted_data_buf[97] : encrypted_data_buf_next[97];   // modexp_top.v(751)
    assign n9567 = rst ? encrypted_data_buf[96] : encrypted_data_buf_next[96];   // modexp_top.v(751)
    assign n9568 = rst ? encrypted_data_buf[95] : encrypted_data_buf_next[95];   // modexp_top.v(751)
    assign n9569 = rst ? encrypted_data_buf[94] : encrypted_data_buf_next[94];   // modexp_top.v(751)
    assign n9570 = rst ? encrypted_data_buf[93] : encrypted_data_buf_next[93];   // modexp_top.v(751)
    assign n9571 = rst ? encrypted_data_buf[92] : encrypted_data_buf_next[92];   // modexp_top.v(751)
    assign n9572 = rst ? encrypted_data_buf[91] : encrypted_data_buf_next[91];   // modexp_top.v(751)
    assign n9573 = rst ? encrypted_data_buf[90] : encrypted_data_buf_next[90];   // modexp_top.v(751)
    assign n9574 = rst ? encrypted_data_buf[89] : encrypted_data_buf_next[89];   // modexp_top.v(751)
    assign n9575 = rst ? encrypted_data_buf[88] : encrypted_data_buf_next[88];   // modexp_top.v(751)
    assign n9576 = rst ? encrypted_data_buf[87] : encrypted_data_buf_next[87];   // modexp_top.v(751)
    assign n9577 = rst ? encrypted_data_buf[86] : encrypted_data_buf_next[86];   // modexp_top.v(751)
    assign n9578 = rst ? encrypted_data_buf[85] : encrypted_data_buf_next[85];   // modexp_top.v(751)
    assign n9579 = rst ? encrypted_data_buf[84] : encrypted_data_buf_next[84];   // modexp_top.v(751)
    assign n9580 = rst ? encrypted_data_buf[83] : encrypted_data_buf_next[83];   // modexp_top.v(751)
    assign n9581 = rst ? encrypted_data_buf[82] : encrypted_data_buf_next[82];   // modexp_top.v(751)
    assign n9582 = rst ? encrypted_data_buf[81] : encrypted_data_buf_next[81];   // modexp_top.v(751)
    assign n9583 = rst ? encrypted_data_buf[80] : encrypted_data_buf_next[80];   // modexp_top.v(751)
    assign n9584 = rst ? encrypted_data_buf[79] : encrypted_data_buf_next[79];   // modexp_top.v(751)
    assign n9585 = rst ? encrypted_data_buf[78] : encrypted_data_buf_next[78];   // modexp_top.v(751)
    assign n9586 = rst ? encrypted_data_buf[77] : encrypted_data_buf_next[77];   // modexp_top.v(751)
    assign n9587 = rst ? encrypted_data_buf[76] : encrypted_data_buf_next[76];   // modexp_top.v(751)
    assign n9588 = rst ? encrypted_data_buf[75] : encrypted_data_buf_next[75];   // modexp_top.v(751)
    assign n9589 = rst ? encrypted_data_buf[74] : encrypted_data_buf_next[74];   // modexp_top.v(751)
    assign n9590 = rst ? encrypted_data_buf[73] : encrypted_data_buf_next[73];   // modexp_top.v(751)
    assign n9591 = rst ? encrypted_data_buf[72] : encrypted_data_buf_next[72];   // modexp_top.v(751)
    assign n9592 = rst ? encrypted_data_buf[71] : encrypted_data_buf_next[71];   // modexp_top.v(751)
    assign n9593 = rst ? encrypted_data_buf[70] : encrypted_data_buf_next[70];   // modexp_top.v(751)
    assign n9594 = rst ? encrypted_data_buf[69] : encrypted_data_buf_next[69];   // modexp_top.v(751)
    assign n9595 = rst ? encrypted_data_buf[68] : encrypted_data_buf_next[68];   // modexp_top.v(751)
    assign n9596 = rst ? encrypted_data_buf[67] : encrypted_data_buf_next[67];   // modexp_top.v(751)
    assign n9597 = rst ? encrypted_data_buf[66] : encrypted_data_buf_next[66];   // modexp_top.v(751)
    assign n9598 = rst ? encrypted_data_buf[65] : encrypted_data_buf_next[65];   // modexp_top.v(751)
    assign n9599 = rst ? encrypted_data_buf[64] : encrypted_data_buf_next[64];   // modexp_top.v(751)
    assign n9600 = rst ? encrypted_data_buf[63] : encrypted_data_buf_next[63];   // modexp_top.v(751)
    assign n9601 = rst ? encrypted_data_buf[62] : encrypted_data_buf_next[62];   // modexp_top.v(751)
    assign n9602 = rst ? encrypted_data_buf[61] : encrypted_data_buf_next[61];   // modexp_top.v(751)
    assign n9603 = rst ? encrypted_data_buf[60] : encrypted_data_buf_next[60];   // modexp_top.v(751)
    assign n9604 = rst ? encrypted_data_buf[59] : encrypted_data_buf_next[59];   // modexp_top.v(751)
    assign n9605 = rst ? encrypted_data_buf[58] : encrypted_data_buf_next[58];   // modexp_top.v(751)
    assign n9606 = rst ? encrypted_data_buf[57] : encrypted_data_buf_next[57];   // modexp_top.v(751)
    assign n9607 = rst ? encrypted_data_buf[56] : encrypted_data_buf_next[56];   // modexp_top.v(751)
    assign n9608 = rst ? encrypted_data_buf[55] : encrypted_data_buf_next[55];   // modexp_top.v(751)
    assign n9609 = rst ? encrypted_data_buf[54] : encrypted_data_buf_next[54];   // modexp_top.v(751)
    assign n9610 = rst ? encrypted_data_buf[53] : encrypted_data_buf_next[53];   // modexp_top.v(751)
    assign n9611 = rst ? encrypted_data_buf[52] : encrypted_data_buf_next[52];   // modexp_top.v(751)
    assign n9612 = rst ? encrypted_data_buf[51] : encrypted_data_buf_next[51];   // modexp_top.v(751)
    assign n9613 = rst ? encrypted_data_buf[50] : encrypted_data_buf_next[50];   // modexp_top.v(751)
    assign n9614 = rst ? encrypted_data_buf[49] : encrypted_data_buf_next[49];   // modexp_top.v(751)
    assign n9615 = rst ? encrypted_data_buf[48] : encrypted_data_buf_next[48];   // modexp_top.v(751)
    assign n9616 = rst ? encrypted_data_buf[47] : encrypted_data_buf_next[47];   // modexp_top.v(751)
    assign n9617 = rst ? encrypted_data_buf[46] : encrypted_data_buf_next[46];   // modexp_top.v(751)
    assign n9618 = rst ? encrypted_data_buf[45] : encrypted_data_buf_next[45];   // modexp_top.v(751)
    assign n9619 = rst ? encrypted_data_buf[44] : encrypted_data_buf_next[44];   // modexp_top.v(751)
    assign n9620 = rst ? encrypted_data_buf[43] : encrypted_data_buf_next[43];   // modexp_top.v(751)
    assign n9621 = rst ? encrypted_data_buf[42] : encrypted_data_buf_next[42];   // modexp_top.v(751)
    assign n9622 = rst ? encrypted_data_buf[41] : encrypted_data_buf_next[41];   // modexp_top.v(751)
    assign n9623 = rst ? encrypted_data_buf[40] : encrypted_data_buf_next[40];   // modexp_top.v(751)
    assign n9624 = rst ? encrypted_data_buf[39] : encrypted_data_buf_next[39];   // modexp_top.v(751)
    assign n9625 = rst ? encrypted_data_buf[38] : encrypted_data_buf_next[38];   // modexp_top.v(751)
    assign n9626 = rst ? encrypted_data_buf[37] : encrypted_data_buf_next[37];   // modexp_top.v(751)
    assign n9627 = rst ? encrypted_data_buf[36] : encrypted_data_buf_next[36];   // modexp_top.v(751)
    assign n9628 = rst ? encrypted_data_buf[35] : encrypted_data_buf_next[35];   // modexp_top.v(751)
    assign n9629 = rst ? encrypted_data_buf[34] : encrypted_data_buf_next[34];   // modexp_top.v(751)
    assign n9630 = rst ? encrypted_data_buf[33] : encrypted_data_buf_next[33];   // modexp_top.v(751)
    assign n9631 = rst ? encrypted_data_buf[32] : encrypted_data_buf_next[32];   // modexp_top.v(751)
    assign n9632 = rst ? encrypted_data_buf[31] : encrypted_data_buf_next[31];   // modexp_top.v(751)
    assign n9633 = rst ? encrypted_data_buf[30] : encrypted_data_buf_next[30];   // modexp_top.v(751)
    assign n9634 = rst ? encrypted_data_buf[29] : encrypted_data_buf_next[29];   // modexp_top.v(751)
    assign n9635 = rst ? encrypted_data_buf[28] : encrypted_data_buf_next[28];   // modexp_top.v(751)
    assign n9636 = rst ? encrypted_data_buf[27] : encrypted_data_buf_next[27];   // modexp_top.v(751)
    assign n9637 = rst ? encrypted_data_buf[26] : encrypted_data_buf_next[26];   // modexp_top.v(751)
    assign n9638 = rst ? encrypted_data_buf[25] : encrypted_data_buf_next[25];   // modexp_top.v(751)
    assign n9639 = rst ? encrypted_data_buf[24] : encrypted_data_buf_next[24];   // modexp_top.v(751)
    assign n9640 = rst ? encrypted_data_buf[23] : encrypted_data_buf_next[23];   // modexp_top.v(751)
    assign n9641 = rst ? encrypted_data_buf[22] : encrypted_data_buf_next[22];   // modexp_top.v(751)
    assign n9642 = rst ? encrypted_data_buf[21] : encrypted_data_buf_next[21];   // modexp_top.v(751)
    assign n9643 = rst ? encrypted_data_buf[20] : encrypted_data_buf_next[20];   // modexp_top.v(751)
    assign n9644 = rst ? encrypted_data_buf[19] : encrypted_data_buf_next[19];   // modexp_top.v(751)
    assign n9645 = rst ? encrypted_data_buf[18] : encrypted_data_buf_next[18];   // modexp_top.v(751)
    assign n9646 = rst ? encrypted_data_buf[17] : encrypted_data_buf_next[17];   // modexp_top.v(751)
    assign n9647 = rst ? encrypted_data_buf[16] : encrypted_data_buf_next[16];   // modexp_top.v(751)
    assign n9648 = rst ? encrypted_data_buf[15] : encrypted_data_buf_next[15];   // modexp_top.v(751)
    assign n9649 = rst ? encrypted_data_buf[14] : encrypted_data_buf_next[14];   // modexp_top.v(751)
    assign n9650 = rst ? encrypted_data_buf[13] : encrypted_data_buf_next[13];   // modexp_top.v(751)
    assign n9651 = rst ? encrypted_data_buf[12] : encrypted_data_buf_next[12];   // modexp_top.v(751)
    assign n9652 = rst ? encrypted_data_buf[11] : encrypted_data_buf_next[11];   // modexp_top.v(751)
    assign n9653 = rst ? encrypted_data_buf[10] : encrypted_data_buf_next[10];   // modexp_top.v(751)
    assign n9654 = rst ? encrypted_data_buf[9] : encrypted_data_buf_next[9];   // modexp_top.v(751)
    assign n9655 = rst ? encrypted_data_buf[8] : encrypted_data_buf_next[8];   // modexp_top.v(751)
    assign n9656 = rst ? encrypted_data_buf[7] : encrypted_data_buf_next[7];   // modexp_top.v(751)
    assign n9657 = rst ? encrypted_data_buf[6] : encrypted_data_buf_next[6];   // modexp_top.v(751)
    assign n9658 = rst ? encrypted_data_buf[5] : encrypted_data_buf_next[5];   // modexp_top.v(751)
    assign n9659 = rst ? encrypted_data_buf[4] : encrypted_data_buf_next[4];   // modexp_top.v(751)
    assign n9660 = rst ? encrypted_data_buf[3] : encrypted_data_buf_next[3];   // modexp_top.v(751)
    assign n9661 = rst ? encrypted_data_buf[2] : encrypted_data_buf_next[2];   // modexp_top.v(751)
    assign n9662 = rst ? encrypted_data_buf[1] : encrypted_data_buf_next[1];   // modexp_top.v(751)
    assign n9663 = rst ? encrypted_data_buf[0] : encrypted_data_buf_next[0];   // modexp_top.v(751)
    VERIFIC_DFFRS i5534 (.d(exp_reg_state_next[1]), .clk(clk), .s(1'b0), 
            .r(rst), .q(exp_state[1]));   // modexp_top.v(751)
    
endmodule

//
// Verific Verilog Description of module reg256byte
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of OPERATOR add_8u_8u
//

module add_8u_8u (cin, a, b, o, cout);
    input cin;
    input [7:0]a;
    input [7:0]b;
    output [7:0]o;
    output cout;
    
    
    wire n2, n4, n6, n8, n10, n12, n14;
    
    VERIFIC_FADD i1 (.cin(cin), .a(a[0]), .b(b[0]), .o(o[0]), .cout(n2));
    VERIFIC_FADD i2 (.cin(n2), .a(a[1]), .b(b[1]), .o(o[1]), .cout(n4));
    VERIFIC_FADD i3 (.cin(n4), .a(a[2]), .b(b[2]), .o(o[2]), .cout(n6));
    VERIFIC_FADD i4 (.cin(n6), .a(a[3]), .b(b[3]), .o(o[3]), .cout(n8));
    VERIFIC_FADD i5 (.cin(n8), .a(a[4]), .b(b[4]), .o(o[4]), .cout(n10));
    VERIFIC_FADD i6 (.cin(n10), .a(a[5]), .b(b[5]), .o(o[5]), .cout(n12));
    VERIFIC_FADD i7 (.cin(n12), .a(a[6]), .b(b[6]), .o(o[6]), .cout(n14));
    VERIFIC_FADD i8 (.cin(n14), .a(a[7]), .b(b[7]), .o(o[7]), .cout(cout));
    
endmodule

//
// Verific Verilog Description of module modexp
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module mem_wr
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module oc8051_xram
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module reg16byte
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module aes_128
// module not written out since it is a black box. 
//

/* verilator coverage_on */
